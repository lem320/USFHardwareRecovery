module rom_error2 (
    input [8:0] address,
    output reg [11:0] data
);

always @(*) begin
    case (address)
        9'h000: data = 12'h7E5;
        9'h001: data = 12'h7E5;
        9'h002: data = 12'h7E5;
        9'h003: data = 12'h7E5;
        9'h004: data = 12'h7E5;
        9'h005: data = 12'h7E5;
        9'h006: data = 12'h7E5;
        9'h007: data = 12'h7E5;
        9'h008: data = 12'h7E5;
        9'h009: data = 12'h7E5;
        9'h00A: data = 12'h7E5;
        9'h00B: data = 12'h7E5;
        9'h00C: data = 12'h7E5;
        9'h00D: data = 12'h7E5;
        9'h00E: data = 12'h7E5;
        9'h00F: data = 12'h7E5;
        9'h010: data = 12'h7E5;
        9'h011: data = 12'h7E5;
        9'h012: data = 12'h7E5;
        9'h013: data = 12'h7E5;
        9'h014: data = 12'h7E5;
        9'h015: data = 12'h7E5;
        9'h016: data = 12'h7E5;
        9'h017: data = 12'h7E5;
        9'h018: data = 12'h7E5;
        9'h019: data = 12'h7E5;
        9'h01A: data = 12'h7E5;
        9'h01B: data = 12'h7E5;
        9'h01C: data = 12'h7E5;
        9'h01D: data = 12'h7E5;
        9'h01E: data = 12'h7E5;
        9'h01F: data = 12'h7E5;
        9'h020: data = 12'h7E5;
        9'h021: data = 12'h7E5;
        9'h022: data = 12'h7E5;
        9'h023: data = 12'h7E5;
        9'h024: data = 12'h7E5;
        9'h025: data = 12'h7E5;
        9'h026: data = 12'h7E5;
        9'h027: data = 12'h7E5;
        9'h028: data = 12'h7E5;
        9'h029: data = 12'h7E5;
        9'h02A: data = 12'h7E5;
        9'h02B: data = 12'h7E5;
        9'h02C: data = 12'h7E5;
        9'h02D: data = 12'h7E5;
        9'h02E: data = 12'h7E5;
        9'h02F: data = 12'h7E5;
        9'h030: data = 12'h7E5;
        9'h031: data = 12'h7E5;
        9'h032: data = 12'h7E5;
        9'h033: data = 12'h7E5;
        9'h034: data = 12'h7E5;
        9'h035: data = 12'h7E5;
        9'h036: data = 12'h7E5;
        9'h037: data = 12'h7E5;
        9'h038: data = 12'h80D;
        9'h039: data = 12'h80D;
        9'h03A: data = 12'h80D;
        9'h03B: data = 12'h80D;
        9'h03C: data = 12'h80D;
        9'h03D: data = 12'h80D;
        9'h03E: data = 12'h80D;
        9'h03F: data = 12'h80D;
        9'h040: data = 12'h80D;
        9'h041: data = 12'h80D;
        9'h042: data = 12'h80D;
        9'h043: data = 12'h80D;
        9'h044: data = 12'h80D;
        9'h045: data = 12'h80D;
        9'h046: data = 12'h80D;
        9'h047: data = 12'h80D;
        9'h048: data = 12'h80D;
        9'h049: data = 12'h80D;
        9'h04A: data = 12'h80D;
        9'h04B: data = 12'h80D;
        9'h04C: data = 12'h80D;
        9'h04D: data = 12'h80D;
        9'h04E: data = 12'h80D;
        9'h04F: data = 12'h80D;
        9'h050: data = 12'h80D;
        9'h051: data = 12'h80D;
        9'h052: data = 12'h80D;
        9'h053: data = 12'h80D;
        9'h054: data = 12'h80D;
        9'h055: data = 12'h80D;
        9'h056: data = 12'h80D;
        9'h057: data = 12'h80A;
        9'h058: data = 12'h80A;
        9'h059: data = 12'h80A;
        9'h05A: data = 12'h80A;
        9'h05B: data = 12'h80A;
        9'h05C: data = 12'h80A;
        9'h05D: data = 12'h80A;
        9'h05E: data = 12'h80A;
        9'h05F: data = 12'h80A;
        9'h060: data = 12'h80A;
        9'h061: data = 12'h80A;
        9'h062: data = 12'h80A;
        9'h063: data = 12'h80A;
        9'h064: data = 12'h80A;
        9'h065: data = 12'h80A;
        9'h066: data = 12'h80A;
        9'h067: data = 12'h80A;
        9'h068: data = 12'h80A;
        9'h069: data = 12'h80A;
        9'h06A: data = 12'h80A;
        9'h06B: data = 12'h80A;
        9'h06C: data = 12'h80A;
        9'h06D: data = 12'h80A;
        9'h06E: data = 12'h80A;
        9'h06F: data = 12'h80A;
        9'h070: data = 12'h80A;
        9'h071: data = 12'h80A;
        9'h072: data = 12'h80A;
        9'h073: data = 12'h80A;
        9'h074: data = 12'h80A;
        9'h075: data = 12'h80A;
        9'h076: data = 12'h28B;
        9'h077: data = 12'h28B;
        9'h078: data = 12'h28B;
        9'h079: data = 12'h28B;
        9'h07A: data = 12'h28B;
        9'h07B: data = 12'h28B;
        9'h07C: data = 12'h28B;
        9'h07D: data = 12'h28B;
        9'h07E: data = 12'h28B;
        9'h07F: data = 12'h28B;
        9'h080: data = 12'h28B;
        9'h081: data = 12'h28B;
        9'h082: data = 12'h28B;
        9'h083: data = 12'h28B;
        9'h084: data = 12'h28B;
        9'h085: data = 12'h28B;
        9'h086: data = 12'h28B;
        9'h087: data = 12'h28B;
        9'h088: data = 12'h28B;
        9'h089: data = 12'h28B;
        9'h08A: data = 12'h28B;
        9'h08B: data = 12'h28B;
        9'h08C: data = 12'h28B;
        9'h08D: data = 12'h28B;
        9'h08E: data = 12'h28B;
        9'h08F: data = 12'h28B;
        9'h090: data = 12'h28B;
        9'h091: data = 12'h28B;
        9'h092: data = 12'h28B;
        9'h093: data = 12'h28B;
        9'h094: data = 12'h28B;
        9'h095: data = 12'h5AA;
        9'h096: data = 12'h5AA;
        9'h097: data = 12'h5AA;
        9'h098: data = 12'h5AA;
        9'h099: data = 12'h5AA;
        9'h09A: data = 12'h5AA;
        9'h09B: data = 12'h5AA;
        9'h09C: data = 12'h5AA;
        9'h09D: data = 12'h5AA;
        9'h09E: data = 12'h5AA;
        9'h09F: data = 12'h5AA;
        9'h0A0: data = 12'h5AA;
        9'h0A1: data = 12'h5AA;
        9'h0A2: data = 12'h5AA;
        9'h0A3: data = 12'h5AA;
        9'h0A4: data = 12'h5AA;
        9'h0A5: data = 12'h5AA;
        9'h0A6: data = 12'h5AA;
        9'h0A7: data = 12'h5AA;
        9'h0A8: data = 12'h5AA;
        9'h0A9: data = 12'h5AA;
        9'h0AA: data = 12'h5AA;
        9'h0AB: data = 12'h5AA;
        9'h0AC: data = 12'h5AA;
        9'h0AD: data = 12'h5AA;
        9'h0AE: data = 12'h5AA;
        9'h0AF: data = 12'h5AA;
        9'h0B0: data = 12'h5AA;
        9'h0B1: data = 12'h5AA;
        9'h0B2: data = 12'h5AA;
        9'h0B3: data = 12'h5AA;
        9'h0B4: data = 12'h7CC;
        9'h0B5: data = 12'h7CC;
        9'h0B6: data = 12'h7CC;
        9'h0B7: data = 12'h7CC;
        9'h0B8: data = 12'h7CC;
        9'h0B9: data = 12'h7CC;
        9'h0BA: data = 12'h7CC;
        9'h0BB: data = 12'h7CC;
        9'h0BC: data = 12'h7CC;
        9'h0BD: data = 12'h7CC;
        9'h0BE: data = 12'h7CC;
        9'h0BF: data = 12'h7CC;
        9'h0C0: data = 12'h7CC;
        9'h0C1: data = 12'h7CC;
        9'h0C2: data = 12'h7CC;
        9'h0C3: data = 12'h7CC;
        9'h0C4: data = 12'h7CC;
        9'h0C5: data = 12'h7CC;
        9'h0C6: data = 12'h7CC;
        9'h0C7: data = 12'h7CC;
        9'h0C8: data = 12'h7CC;
        9'h0C9: data = 12'h7CC;
        9'h0CA: data = 12'h7CC;
        9'h0CB: data = 12'h7CC;
        9'h0CC: data = 12'h7CC;
        9'h0CD: data = 12'h7CC;
        9'h0CE: data = 12'h7CC;
        9'h0CF: data = 12'h7CC;
        9'h0D0: data = 12'h7CC;
        9'h0D1: data = 12'h7CC;
        9'h0D2: data = 12'h7CC;
        9'h0D3: data = 12'h066;
        9'h0D4: data = 12'h066;
        9'h0D5: data = 12'h066;
        9'h0D6: data = 12'h066;
        9'h0D7: data = 12'h066;
        9'h0D8: data = 12'h066;
        9'h0D9: data = 12'h066;
        9'h0DA: data = 12'h066;
        9'h0DB: data = 12'h066;
        9'h0DC: data = 12'h066;
        9'h0DD: data = 12'h066;
        9'h0DE: data = 12'h066;
        9'h0DF: data = 12'h066;
        9'h0E0: data = 12'h066;
        9'h0E1: data = 12'h066;
        9'h0E2: data = 12'h066;
        9'h0E3: data = 12'h066;
        9'h0E4: data = 12'h066;
        9'h0E5: data = 12'h066;
        9'h0E6: data = 12'h066;
        9'h0E7: data = 12'h066;
        9'h0E8: data = 12'h066;
        9'h0E9: data = 12'h066;
        9'h0EA: data = 12'h066;
        9'h0EB: data = 12'h066;
        9'h0EC: data = 12'h066;
        9'h0ED: data = 12'h066;
        9'h0EE: data = 12'h066;
        9'h0EF: data = 12'h066;
        9'h0F0: data = 12'h066;
        9'h0F1: data = 12'h066;
        9'h0F2: data = 12'h05B;
        9'h0F3: data = 12'h05B;
        9'h0F4: data = 12'h05B;
        9'h0F5: data = 12'h05B;
        9'h0F6: data = 12'h05B;
        9'h0F7: data = 12'h05B;
        9'h0F8: data = 12'h05B;
        9'h0F9: data = 12'h05B;
        9'h0FA: data = 12'h05B;
        9'h0FB: data = 12'h05B;
        9'h0FC: data = 12'h05B;
        9'h0FD: data = 12'h05B;
        9'h0FE: data = 12'h05B;
        9'h0FF: data = 12'h05B;
        9'h100: data = 12'h05B;
        9'h101: data = 12'h05B;
        9'h102: data = 12'h05B;
        9'h103: data = 12'h05B;
        9'h104: data = 12'h05B;
        9'h105: data = 12'h05B;
        9'h106: data = 12'h05B;
        9'h107: data = 12'h05B;
        9'h108: data = 12'h05B;
        9'h109: data = 12'h05B;
        9'h10A: data = 12'h05B;
        9'h10B: data = 12'h05B;
        9'h10C: data = 12'h05B;
        9'h10D: data = 12'h05B;
        9'h10E: data = 12'h05B;
        9'h10F: data = 12'h05B;
        9'h110: data = 12'h05B;
        9'h111: data = 12'h07E;
        9'h112: data = 12'h07E;
        9'h113: data = 12'h07E;
        9'h114: data = 12'h07E;
        9'h115: data = 12'h07E;
        9'h116: data = 12'h07E;
        9'h117: data = 12'h07E;
        9'h118: data = 12'h07E;
        9'h119: data = 12'h07E;
        9'h11A: data = 12'h07E;
        9'h11B: data = 12'h07E;
        9'h11C: data = 12'h07E;
        9'h11D: data = 12'h07E;
        9'h11E: data = 12'h07E;
        9'h11F: data = 12'h07E;
        9'h120: data = 12'h07E;
        9'h121: data = 12'h07E;
        9'h122: data = 12'h07E;
        9'h123: data = 12'h07E;
        9'h124: data = 12'h07E;
        9'h125: data = 12'h07E;
        9'h126: data = 12'h07E;
        9'h127: data = 12'h07E;
        9'h128: data = 12'h07E;
        9'h129: data = 12'h07E;
        9'h12A: data = 12'h07E;
        9'h12B: data = 12'h07E;
        9'h12C: data = 12'h07E;
        9'h12D: data = 12'h07E;
        9'h12E: data = 12'h07E;
        9'h12F: data = 12'h07E;
        9'h130: data = 12'h07F;
        9'h131: data = 12'h07F;
        9'h132: data = 12'h07F;
        9'h133: data = 12'h07F;
        9'h134: data = 12'h07F;
        9'h135: data = 12'h07F;
        9'h136: data = 12'h07F;
        9'h137: data = 12'h07F;
        9'h138: data = 12'h07F;
        9'h139: data = 12'h07F;
        9'h13A: data = 12'h07F;
        9'h13B: data = 12'h07F;
        9'h13C: data = 12'h07F;
        9'h13D: data = 12'h07F;
        9'h13E: data = 12'h07F;
        9'h13F: data = 12'h07F;
        9'h140: data = 12'h07F;
        9'h141: data = 12'h07F;
        9'h142: data = 12'h07F;
        9'h143: data = 12'h07F;
        9'h144: data = 12'h07F;
        9'h145: data = 12'h07F;
        9'h146: data = 12'h07F;
        9'h147: data = 12'h07F;
        9'h148: data = 12'h07F;
        9'h149: data = 12'h07F;
        9'h14A: data = 12'h07F;
        9'h14B: data = 12'h07F;
        9'h14C: data = 12'h07F;
        9'h14D: data = 12'h07F;
        9'h14E: data = 12'h07F;
        9'h14F: data = 12'h08B;
        9'h150: data = 12'h08B;
        9'h151: data = 12'h08B;
        9'h152: data = 12'h08B;
        9'h153: data = 12'h08B;
        9'h154: data = 12'h08B;
        9'h155: data = 12'h08B;
        9'h156: data = 12'h08B;
        9'h157: data = 12'h08B;
        9'h158: data = 12'h08B;
        9'h159: data = 12'h08B;
        9'h15A: data = 12'h08B;
        9'h15B: data = 12'h08B;
        9'h15C: data = 12'h08B;
        9'h15D: data = 12'h08B;
        9'h15E: data = 12'h08B;
        9'h15F: data = 12'h08B;
        9'h160: data = 12'h08B;
        9'h161: data = 12'h08B;
        9'h162: data = 12'h08B;
        9'h163: data = 12'h08B;
        9'h164: data = 12'h08B;
        9'h165: data = 12'h08B;
        9'h166: data = 12'h08B;
        9'h167: data = 12'h08B;
        9'h168: data = 12'h08B;
        9'h169: data = 12'h08B;
        9'h16A: data = 12'h08B;
        9'h16B: data = 12'h08B;
        9'h16C: data = 12'h08B;
        9'h16D: data = 12'h08B;
        9'h16E: data = 12'h0A2;
        9'h16F: data = 12'h0A2;
        9'h170: data = 12'h0A2;
        9'h171: data = 12'h0A2;
        9'h172: data = 12'h0A2;
        9'h173: data = 12'h0A2;
        9'h174: data = 12'h0A2;
        9'h175: data = 12'h0A2;
        9'h176: data = 12'h0A2;
        9'h177: data = 12'h0A2;
        9'h178: data = 12'h0A2;
        9'h179: data = 12'h0A2;
        9'h17A: data = 12'h0A2;
        9'h17B: data = 12'h0A2;
        9'h17C: data = 12'h0A2;
        9'h17D: data = 12'h0A2;
        9'h17E: data = 12'h0A2;
        9'h17F: data = 12'h0A2;
        9'h180: data = 12'h0A2;
        9'h181: data = 12'h0A2;
        9'h182: data = 12'h0A2;
        9'h183: data = 12'h0A2;
        9'h184: data = 12'h0A2;
        9'h185: data = 12'h0A2;
        9'h186: data = 12'h0A2;
        9'h187: data = 12'h0A2;
        9'h188: data = 12'h0A2;
        9'h189: data = 12'h0A2;
        9'h18A: data = 12'h0A2;
        9'h18B: data = 12'h0A2;
        9'h18C: data = 12'h0A2;
        9'h18D: data = 12'h0A5;
        9'h18E: data = 12'h0A5;
        9'h18F: data = 12'h0A5;
        9'h190: data = 12'h0A5;
        9'h191: data = 12'h0A5;
        9'h192: data = 12'h0A5;
        9'h193: data = 12'h0A5;
        9'h194: data = 12'h0A5;
        9'h195: data = 12'h0A5;
        9'h196: data = 12'h0A5;
        9'h197: data = 12'h0A5;
        9'h198: data = 12'h0A5;
        9'h199: data = 12'h0A5;
        9'h19A: data = 12'h0A5;
        9'h19B: data = 12'h0A5;
        9'h19C: data = 12'h0A5;
        9'h19D: data = 12'h0A5;
        9'h19E: data = 12'h0A5;
        9'h19F: data = 12'h0A5;
        9'h1A0: data = 12'h0A5;
        9'h1A1: data = 12'h0A5;
        9'h1A2: data = 12'h0A5;
        9'h1A3: data = 12'h0A5;
        9'h1A4: data = 12'h0A5;
        9'h1A5: data = 12'h0A5;
        9'h1A6: data = 12'h0A5;
        9'h1A7: data = 12'h0A5;
        9'h1A8: data = 12'h0A5;
        9'h1A9: data = 12'h0A5;
        9'h1AA: data = 12'h0A5;
        9'h1AB: data = 12'h0A5;
        9'h1AC: data = 12'h0BC;
        9'h1AD: data = 12'h0BC;
        9'h1AE: data = 12'h0BC;
        9'h1AF: data = 12'h0BC;
        9'h1B0: data = 12'h0BC;
        9'h1B1: data = 12'h0BC;
        9'h1B2: data = 12'h0BC;
        9'h1B3: data = 12'h0BC;
        9'h1B4: data = 12'h0BC;
        9'h1B5: data = 12'h0BC;
        9'h1B6: data = 12'h0BC;
        9'h1B7: data = 12'h0BC;
        9'h1B8: data = 12'h0BC;
        9'h1B9: data = 12'h0BC;
        9'h1BA: data = 12'h0BC;
        9'h1BB: data = 12'h0BC;
        9'h1BC: data = 12'h0BC;
        9'h1BD: data = 12'h0BC;
        9'h1BE: data = 12'h0BC;
        9'h1BF: data = 12'h0BC;
        9'h1C0: data = 12'h0BC;
        9'h1C1: data = 12'h0BC;
        9'h1C2: data = 12'h0BC;
        9'h1C3: data = 12'h0BC;
        9'h1C4: data = 12'h0BC;
        9'h1C5: data = 12'h0BC;
        9'h1C6: data = 12'h0BC;
        9'h1C7: data = 12'h0BC;
        9'h1C8: data = 12'h0BC;
        9'h1C9: data = 12'h0BC;
        9'h1CA: data = 12'h0BC;
        9'h1CB: data = 12'h0C9;
        9'h1CC: data = 12'h0C9;
        9'h1CD: data = 12'h0C9;
        9'h1CE: data = 12'h0C9;
        9'h1CF: data = 12'h0C9;
        9'h1D0: data = 12'h0C9;
        9'h1D1: data = 12'h0C9;
        9'h1D2: data = 12'h0C9;
        9'h1D3: data = 12'h0C9;
        9'h1D4: data = 12'h0C9;
        9'h1D5: data = 12'h0C9;
        9'h1D6: data = 12'h0C9;
        9'h1D7: data = 12'h0C9;
        9'h1D8: data = 12'h0C9;
        9'h1D9: data = 12'h0C9;
        9'h1DA: data = 12'h0C9;
        9'h1DB: data = 12'h0C9;
        9'h1DC: data = 12'h0C9;
        9'h1DD: data = 12'h0C9;
        9'h1DE: data = 12'h0C9;
        9'h1DF: data = 12'h0C9;
        9'h1E0: data = 12'h0C9;
        9'h1E1: data = 12'h0C9;
        9'h1E2: data = 12'h0C9;
        9'h1E3: data = 12'h0C9;
        9'h1E4: data = 12'h0C9;
        9'h1E5: data = 12'h0C9;
        9'h1E6: data = 12'h0C9;
        9'h1E7: data = 12'h0C9;
        9'h1E8: data = 12'h0C9;
        9'h1E9: data = 12'h0C9;
        9'h1EA: data = 12'h0E5;
        9'h1EB: data = 12'h0E5;
        9'h1EC: data = 12'h0E5;
        9'h1ED: data = 12'h0E5;
        9'h1EE: data = 12'h0E5;
        9'h1EF: data = 12'h0E5;
        9'h1F0: data = 12'h0E5;
        9'h1F1: data = 12'h0E5;
        9'h1F2: data = 12'h0E5;
        9'h1F3: data = 12'h0E5;
        9'h1F4: data = 12'h0E5;
        9'h1F5: data = 12'h0E5;
        9'h1F6: data = 12'h0E5;
        9'h1F7: data = 12'h0E5;
        9'h1F8: data = 12'h0E5;
        9'h1F9: data = 12'h0E5;
        9'h1FA: data = 12'h0E5;
        9'h1FB: data = 12'h0E5;
        9'h1FC: data = 12'h0E5;
        9'h1FD: data = 12'h0E5;
        9'h1FE: data = 12'h0E5;
        9'h1FF: data = 12'h0E5;
        default: data = 12'h000;
    endcase
end

endmodule

module rom_test1 (
    input [14:0] address,
    output reg [11:0] data
);

always @(*) begin
    case (address)
        15'h0000: data = 12'h78F;
        15'h0001: data = 12'h790;
        15'h0002: data = 12'h79F;
        15'h0003: data = 12'h7A6;
        15'h0004: data = 12'h7AD;
        15'h0005: data = 12'h7B9;
        15'h0006: data = 12'h7C3;
        15'h0007: data = 12'h7D2;
        15'h0008: data = 12'h7D9;
        15'h0009: data = 12'h7E3;
        15'h000A: data = 12'h7E7;
        15'h000B: data = 12'h7F1;
        15'h000C: data = 12'h7F3;
        15'h000D: data = 12'h7FB;
        15'h000E: data = 12'h806;
        15'h000F: data = 12'h80C;
        15'h0010: data = 12'h812;
        15'h0011: data = 12'h815;
        15'h0012: data = 12'h095;
        15'h0013: data = 12'h0A0;
        15'h0014: data = 12'h70B;
        15'h0015: data = 12'h71C;
        15'h0016: data = 12'h725;
        15'h0017: data = 12'h72D;
        15'h0018: data = 12'h735;
        15'h0019: data = 12'h744;
        15'h001A: data = 12'h74D;
        15'h001B: data = 12'h75C;
        15'h001C: data = 12'h765;
        15'h001D: data = 12'h778;
        15'h001E: data = 12'h782;
        15'h001F: data = 12'h78F;
        15'h0020: data = 12'h7B5;
        15'h0021: data = 12'h0C5;
        15'h0022: data = 12'h7C6;
        15'h0023: data = 12'h7CA;
        15'h0024: data = 12'h7D5;
        15'h0025: data = 12'h7DC;
        15'h0026: data = 12'h7E4;
        15'h0027: data = 12'h7F0;
        15'h0028: data = 12'h7F8;
        15'h0029: data = 12'h7F5;
        15'h002A: data = 12'h801;
        15'h002B: data = 12'h805;
        15'h002C: data = 12'h2E9;
        15'h002D: data = 12'h088;
        15'h002E: data = 12'h095;
        15'h002F: data = 12'h09A;
        15'h0030: data = 12'h09C;
        15'h0031: data = 12'h0AA;
        15'h0032: data = 12'h0AD;
        15'h0033: data = 12'h0BA;
        15'h0034: data = 12'h0BB;
        15'h0035: data = 12'h0BB;
        15'h0036: data = 12'h0C6;
        15'h0037: data = 12'h0C8;
        15'h0038: data = 12'h0C9;
        15'h0039: data = 12'h0CB;
        15'h003A: data = 12'h0D4;
        15'h003B: data = 12'h0D3;
        15'h003C: data = 12'h0D1;
        15'h003D: data = 12'h0CE;
        15'h003E: data = 12'h0CF;
        15'h003F: data = 12'h0CA;
        15'h0040: data = 12'h0C5;
        15'h0041: data = 12'h0BE;
        15'h0042: data = 12'h0B9;
        15'h0043: data = 12'h0BA;
        15'h0044: data = 12'h0BC;
        15'h0045: data = 12'h0BD;
        15'h0046: data = 12'h0B9;
        15'h0047: data = 12'h0BD;
        15'h0048: data = 12'h0BB;
        15'h0049: data = 12'h0BE;
        15'h004A: data = 12'h0BB;
        15'h004B: data = 12'h0B8;
        15'h004C: data = 12'h0B1;
        15'h004D: data = 12'h0AE;
        15'h004E: data = 12'h0A4;
        15'h004F: data = 12'h09A;
        15'h0050: data = 12'h095;
        15'h0051: data = 12'h08A;
        15'h0052: data = 12'h082;
        15'h0053: data = 12'h082;
        15'h0054: data = 12'h07F;
        15'h0055: data = 12'h084;
        15'h0056: data = 12'h07F;
        15'h0057: data = 12'h078;
        15'h0058: data = 12'h06F;
        15'h0059: data = 12'h063;
        15'h005A: data = 12'h053;
        15'h005B: data = 12'h046;
        15'h005C: data = 12'h040;
        15'h005D: data = 12'h017;
        15'h005E: data = 12'h7BF;
        15'h005F: data = 12'h7B7;
        15'h0060: data = 12'h7B0;
        15'h0061: data = 12'h7A9;
        15'h0062: data = 12'h793;
        15'h0063: data = 12'h782;
        15'h0064: data = 12'h768;
        15'h0065: data = 12'h760;
        15'h0066: data = 12'h751;
        15'h0067: data = 12'h74B;
        15'h0068: data = 12'h745;
        15'h0069: data = 12'h740;
        15'h006A: data = 12'h735;
        15'h006B: data = 12'h728;
        15'h006C: data = 12'h717;
        15'h006D: data = 12'h700;
        15'h006E: data = 12'h6E9;
        15'h006F: data = 12'h6D6;
        15'h0070: data = 12'h6D0;
        15'h0071: data = 12'h6C7;
        15'h0072: data = 12'h6BE;
        15'h0073: data = 12'h6B5;
        15'h0074: data = 12'h6A5;
        15'h0075: data = 12'h698;
        15'h0076: data = 12'h686;
        15'h0077: data = 12'h674;
        15'h0078: data = 12'h665;
        15'h0079: data = 12'h64A;
        15'h007A: data = 12'h637;
        15'h007B: data = 12'h626;
        15'h007C: data = 12'h619;
        15'h007D: data = 12'h607;
        15'h007E: data = 12'h5F9;
        15'h007F: data = 12'h5EF;
        15'h0080: data = 12'h5E0;
        15'h0081: data = 12'h5CC;
        15'h0082: data = 12'h5C4;
        15'h0083: data = 12'h5B2;
        15'h0084: data = 12'h59E;
        15'h0085: data = 12'h589;
        15'h0086: data = 12'h570;
        15'h0087: data = 12'h560;
        15'h0088: data = 12'h54B;
        15'h0089: data = 12'h532;
        15'h008A: data = 12'h519;
        15'h008B: data = 12'h50B;
        15'h008C: data = 12'h4F7;
        15'h008D: data = 12'h4E4;
        15'h008E: data = 12'h4CD;
        15'h008F: data = 12'h4C0;
        15'h0090: data = 12'h4AE;
        15'h0091: data = 12'h49D;
        15'h0092: data = 12'h48B;
        15'h0093: data = 12'h478;
        15'h0094: data = 12'h461;
        15'h0095: data = 12'h455;
        15'h0096: data = 12'h43D;
        15'h0097: data = 12'h429;
        15'h0098: data = 12'h411;
        15'h0099: data = 12'h3FE;
        15'h009A: data = 12'h3E9;
        15'h009B: data = 12'h3D4;
        15'h009C: data = 12'h3BA;
        15'h009D: data = 12'h3A1;
        15'h009E: data = 12'h38E;
        15'h009F: data = 12'h373;
        15'h00A0: data = 12'h35F;
        15'h00A1: data = 12'h346;
        15'h00A2: data = 12'h334;
        15'h00A3: data = 12'h31A;
        15'h00A4: data = 12'h301;
        15'h00A5: data = 12'h2EC;
        15'h00A6: data = 12'h2D4;
        15'h00A7: data = 12'h2BB;
        15'h00A8: data = 12'h2A5;
        15'h00A9: data = 12'h28A;
        15'h00AA: data = 12'h277;
        15'h00AB: data = 12'h25F;
        15'h00AC: data = 12'h244;
        15'h00AD: data = 12'h232;
        15'h00AE: data = 12'h210;
        15'h00AF: data = 12'h1FB;
        15'h00B0: data = 12'h1E7;
        15'h00B1: data = 12'h1CE;
        15'h00B2: data = 12'h1B1;
        15'h00B3: data = 12'h19C;
        15'h00B4: data = 12'h184;
        15'h00B5: data = 12'h16B;
        15'h00B6: data = 12'h151;
        15'h00B7: data = 12'h140;
        15'h00B8: data = 12'h126;
        15'h00B9: data = 12'h10F;
        15'h00BA: data = 12'h0F7;
        15'h00BB: data = 12'h0DF;
        15'h00BC: data = 12'h0CA;
        15'h00BD: data = 12'h0B0;
        15'h00BE: data = 12'h097;
        15'h00BF: data = 12'h084;
        15'h00C0: data = 12'h06E;
        15'h00C1: data = 12'h057;
        15'h00C2: data = 12'h03A;
        15'h00C3: data = 12'h7A8;
        15'h00C4: data = 12'h7C0;
        15'h00C5: data = 12'h7A9;
        15'h00C6: data = 12'h790;
        15'h00C7: data = 12'h779;
        15'h00C8: data = 12'h763;
        15'h00C9: data = 12'h74C;
        15'h00CA: data = 12'h738;
        15'h00CB: data = 12'h723;
        15'h00CC: data = 12'h70D;
        15'h00CD: data = 12'h6F7;
        15'h00CE: data = 12'h6DD;
        15'h00CF: data = 12'h6C6;
        15'h00D0: data = 12'h6B3;
        15'h00D1: data = 12'h69B;
        15'h00D2: data = 12'h689;
        15'h00D3: data = 12'h676;
        15'h00D4: data = 12'h65C;
        15'h00D5: data = 12'h649;
        15'h00D6: data = 12'h633;
        15'h00D7: data = 12'h61C;
        15'h00D8: data = 12'h607;
        15'h00D9: data = 12'h5F1;
        15'h00DA: data = 12'h5D9;
        15'h00DB: data = 12'h5C3;
        15'h00DC: data = 12'h5B7;
        15'h00DD: data = 12'h59E;
        15'h00DE: data = 12'h589;
        15'h00DF: data = 12'h579;
        15'h00E0: data = 12'h564;
        15'h00E1: data = 12'h555;
        15'h00E2: data = 12'h541;
        15'h00E3: data = 12'h52B;
        15'h00E4: data = 12'h518;
        15'h00E5: data = 12'h505;
        15'h00E6: data = 12'h4F2;
        15'h00E7: data = 12'h4E0;
        15'h00E8: data = 12'h4C8;
        15'h00E9: data = 12'h4B7;
        15'h00EA: data = 12'h4A0;
        15'h00EB: data = 12'h491;
        15'h00EC: data = 12'h479;
        15'h00ED: data = 12'h463;
        15'h00EE: data = 12'h454;
        15'h00EF: data = 12'h442;
        15'h00F0: data = 12'h426;
        15'h00F1: data = 12'h417;
        15'h00F2: data = 12'h3FF;
        15'h00F3: data = 12'h3EC;
        15'h00F4: data = 12'h3D8;
        15'h00F5: data = 12'h3C5;
        15'h00F6: data = 12'h3AC;
        15'h00F7: data = 12'h39F;
        15'h00F8: data = 12'h390;
        15'h00F9: data = 12'h383;
        15'h00FA: data = 12'h373;
        15'h00FB: data = 12'h361;
        15'h00FC: data = 12'h352;
        15'h00FD: data = 12'h346;
        15'h00FE: data = 12'h33A;
        15'h00FF: data = 12'h330;
        15'h0100: data = 12'h322;
        15'h0101: data = 12'h30E;
        15'h0102: data = 12'h302;
        15'h0103: data = 12'h2F4;
        15'h0104: data = 12'h2E3;
        15'h0105: data = 12'h2D9;
        15'h0106: data = 12'h2C5;
        15'h0107: data = 12'h2B3;
        15'h0108: data = 12'h2A0;
        15'h0109: data = 12'h291;
        15'h010A: data = 12'h280;
        15'h010B: data = 12'h271;
        15'h010C: data = 12'h268;
        15'h010D: data = 12'h25D;
        15'h010E: data = 12'h257;
        15'h010F: data = 12'h249;
        15'h0110: data = 12'h247;
        15'h0111: data = 12'h238;
        15'h0112: data = 12'h238;
        15'h0113: data = 12'h226;
        15'h0114: data = 12'h223;
        15'h0115: data = 12'h217;
        15'h0116: data = 12'h210;
        15'h0117: data = 12'h1FF;
        15'h0118: data = 12'h1F1;
        15'h0119: data = 12'h1E6;
        15'h011A: data = 12'h1D9;
        15'h011B: data = 12'h1D1;
        15'h011C: data = 12'h1C5;
        15'h011D: data = 12'h1BE;
        15'h011E: data = 12'h1BB;
        15'h011F: data = 12'h1B8;
        15'h0120: data = 12'h1B2;
        15'h0121: data = 12'h1B1;
        15'h0122: data = 12'h1A9;
        15'h0123: data = 12'h1A8;
        15'h0124: data = 12'h1A6;
        15'h0125: data = 12'h19A;
        15'h0126: data = 12'h193;
        15'h0127: data = 12'h191;
        15'h0128: data = 12'h185;
        15'h0129: data = 12'h17B;
        15'h012A: data = 12'h177;
        15'h012B: data = 12'h16F;
        15'h012C: data = 12'h16A;
        15'h012D: data = 12'h163;
        15'h012E: data = 12'h168;
        15'h012F: data = 12'h169;
        15'h0130: data = 12'h165;
        15'h0131: data = 12'h16D;
        15'h0132: data = 12'h16E;
        15'h0133: data = 12'h170;
        15'h0134: data = 12'h164;
        15'h0135: data = 12'h165;
        15'h0136: data = 12'h168;
        15'h0137: data = 12'h163;
        15'h0138: data = 12'h15E;
        15'h0139: data = 12'h15C;
        15'h013A: data = 12'h158;
        15'h013B: data = 12'h158;
        15'h013C: data = 12'h15D;
        15'h013D: data = 12'h15D;
        15'h013E: data = 12'h162;
        15'h013F: data = 12'h165;
        15'h0140: data = 12'h16F;
        15'h0141: data = 12'h174;
        15'h0142: data = 12'h177;
        15'h0143: data = 12'h17E;
        15'h0144: data = 12'h180;
        15'h0145: data = 12'h183;
        15'h0146: data = 12'h189;
        15'h0147: data = 12'h18A;
        15'h0148: data = 12'h18F;
        15'h0149: data = 12'h18A;
        15'h014A: data = 12'h18E;
        15'h014B: data = 12'h192;
        15'h014C: data = 12'h19A;
        15'h014D: data = 12'h19C;
        15'h014E: data = 12'h1A1;
        15'h014F: data = 12'h1AD;
        15'h0150: data = 12'h1B6;
        15'h0151: data = 12'h1C4;
        15'h0152: data = 12'h1CF;
        15'h0153: data = 12'h1D9;
        15'h0154: data = 12'h1DE;
        15'h0155: data = 12'h1E9;
        15'h0156: data = 12'h1F2;
        15'h0157: data = 12'h1F7;
        15'h0158: data = 12'h206;
        15'h0159: data = 12'h20A;
        15'h015A: data = 12'h210;
        15'h015B: data = 12'h20F;
        15'h015C: data = 12'h21F;
        15'h015D: data = 12'h225;
        15'h015E: data = 12'h232;
        15'h015F: data = 12'h23C;
        15'h0160: data = 12'h249;
        15'h0161: data = 12'h258;
        15'h0162: data = 12'h267;
        15'h0163: data = 12'h277;
        15'h0164: data = 12'h288;
        15'h0165: data = 12'h293;
        15'h0166: data = 12'h2A4;
        15'h0167: data = 12'h2B3;
        15'h0168: data = 12'h2C1;
        15'h0169: data = 12'h2CD;
        15'h016A: data = 12'h2DD;
        15'h016B: data = 12'h2E7;
        15'h016C: data = 12'h2F6;
        15'h016D: data = 12'h2FE;
        15'h016E: data = 12'h30B;
        15'h016F: data = 12'h319;
        15'h0170: data = 12'h322;
        15'h0171: data = 12'h32E;
        15'h0172: data = 12'h341;
        15'h0173: data = 12'h352;
        15'h0174: data = 12'h365;
        15'h0175: data = 12'h37A;
        15'h0176: data = 12'h390;
        15'h0177: data = 12'h39E;
        15'h0178: data = 12'h3B7;
        15'h0179: data = 12'h3C4;
        15'h017A: data = 12'h3D8;
        15'h017B: data = 12'h3F0;
        15'h017C: data = 12'h403;
        15'h017D: data = 12'h410;
        15'h017E: data = 12'h421;
        15'h017F: data = 12'h435;
        15'h0180: data = 12'h43E;
        15'h0181: data = 12'h456;
        15'h0182: data = 12'h45E;
        15'h0183: data = 12'h472;
        15'h0184: data = 12'h484;
        15'h0185: data = 12'h497;
        15'h0186: data = 12'h4A4;
        15'h0187: data = 12'h4C1;
        15'h0188: data = 12'h4CF;
        15'h0189: data = 12'h4E3;
        15'h018A: data = 12'h4FD;
        15'h018B: data = 12'h513;
        15'h018C: data = 12'h52C;
        15'h018D: data = 12'h543;
        15'h018E: data = 12'h55D;
        15'h018F: data = 12'h573;
        15'h0190: data = 12'h587;
        15'h0191: data = 12'h59D;
        15'h0192: data = 12'h5AE;
        15'h0193: data = 12'h5C1;
        15'h0194: data = 12'h5DC;
        15'h0195: data = 12'h5F0;
        15'h0196: data = 12'h603;
        15'h0197: data = 12'h61A;
        15'h0198: data = 12'h625;
        15'h0199: data = 12'h637;
        15'h019A: data = 12'h64F;
        15'h019B: data = 12'h661;
        15'h019C: data = 12'h679;
        15'h019D: data = 12'h68F;
        15'h019E: data = 12'h6A8;
        15'h019F: data = 12'h6BF;
        15'h01A0: data = 12'h6D5;
        15'h01A1: data = 12'h6ED;
        15'h01A2: data = 12'h708;
        15'h01A3: data = 12'h724;
        15'h01A4: data = 12'h73C;
        15'h01A5: data = 12'h752;
        15'h01A6: data = 12'h76A;
        15'h01A7: data = 12'h783;
        15'h01A8: data = 12'h79D;
        15'h01A9: data = 12'h7B3;
        15'h01AA: data = 12'h7CA;
        15'h01AB: data = 12'h7DC;
        15'h01AC: data = 12'h7F1;
        15'h01AD: data = 12'h80A;
        15'h01AE: data = 12'h06D;
        15'h01AF: data = 12'h085;
        15'h01B0: data = 12'h098;
        15'h01B1: data = 12'h0A8;
        15'h01B2: data = 12'h0BD;
        15'h01B3: data = 12'h0D5;
        15'h01B4: data = 12'h0EE;
        15'h01B5: data = 12'h0FB;
        15'h01B6: data = 12'h118;
        15'h01B7: data = 12'h131;
        15'h01B8: data = 12'h149;
        15'h01B9: data = 12'h161;
        15'h01BA: data = 12'h17C;
        15'h01BB: data = 12'h195;
        15'h01BC: data = 12'h1B0;
        15'h01BD: data = 12'h1C6;
        15'h01BE: data = 12'h1DE;
        15'h01BF: data = 12'h1FC;
        15'h01C0: data = 12'h217;
        15'h01C1: data = 12'h228;
        15'h01C2: data = 12'h240;
        15'h01C3: data = 12'h25B;
        15'h01C4: data = 12'h26F;
        15'h01C5: data = 12'h280;
        15'h01C6: data = 12'h298;
        15'h01C7: data = 12'h2B4;
        15'h01C8: data = 12'h2CD;
        15'h01C9: data = 12'h2DA;
        15'h01CA: data = 12'h2F1;
        15'h01CB: data = 12'h303;
        15'h01CC: data = 12'h31F;
        15'h01CD: data = 12'h32C;
        15'h01CE: data = 12'h343;
        15'h01CF: data = 12'h358;
        15'h01D0: data = 12'h36E;
        15'h01D1: data = 12'h385;
        15'h01D2: data = 12'h397;
        15'h01D3: data = 12'h3B0;
        15'h01D4: data = 12'h3C6;
        15'h01D5: data = 12'h3DC;
        15'h01D6: data = 12'h3F0;
        15'h01D7: data = 12'h405;
        15'h01D8: data = 12'h41E;
        15'h01D9: data = 12'h434;
        15'h01DA: data = 12'h446;
        15'h01DB: data = 12'h45C;
        15'h01DC: data = 12'h474;
        15'h01DD: data = 12'h48F;
        15'h01DE: data = 12'h4A3;
        15'h01DF: data = 12'h4B8;
        15'h01E0: data = 12'h4CB;
        15'h01E1: data = 12'h4E1;
        15'h01E2: data = 12'h4F8;
        15'h01E3: data = 12'h50E;
        15'h01E4: data = 12'h519;
        15'h01E5: data = 12'h532;
        15'h01E6: data = 12'h54C;
        15'h01E7: data = 12'h559;
        15'h01E8: data = 12'h56E;
        15'h01E9: data = 12'h57F;
        15'h01EA: data = 12'h592;
        15'h01EB: data = 12'h5A4;
        15'h01EC: data = 12'h5B5;
        15'h01ED: data = 12'h5C9;
        15'h01EE: data = 12'h5D4;
        15'h01EF: data = 12'h5E8;
        15'h01F0: data = 12'h5F9;
        15'h01F1: data = 12'h610;
        15'h01F2: data = 12'h61D;
        15'h01F3: data = 12'h629;
        15'h01F4: data = 12'h638;
        15'h01F5: data = 12'h641;
        15'h01F6: data = 12'h652;
        15'h01F7: data = 12'h667;
        15'h01F8: data = 12'h675;
        15'h01F9: data = 12'h682;
        15'h01FA: data = 12'h692;
        15'h01FB: data = 12'h69D;
        15'h01FC: data = 12'h6A6;
        15'h01FD: data = 12'h6B9;
        15'h01FE: data = 12'h6C7;
        15'h01FF: data = 12'h6D0;
        15'h0200: data = 12'h6DF;
        15'h0201: data = 12'h6ED;
        15'h0202: data = 12'h6F8;
        15'h0203: data = 12'h703;
        15'h0204: data = 12'h714;
        15'h0205: data = 12'h71E;
        15'h0206: data = 12'h726;
        15'h0207: data = 12'h72C;
        15'h0208: data = 12'h73D;
        15'h0209: data = 12'h74C;
        15'h020A: data = 12'h755;
        15'h020B: data = 12'h764;
        15'h020C: data = 12'h76A;
        15'h020D: data = 12'h77C;
        15'h020E: data = 12'h787;
        15'h020F: data = 12'h78D;
        15'h0210: data = 12'h794;
        15'h0211: data = 12'h79F;
        15'h0212: data = 12'h7A9;
        15'h0213: data = 12'h7B5;
        15'h0214: data = 12'h7BF;
        15'h0215: data = 12'h7C5;
        15'h0216: data = 12'h7CE;
        15'h0217: data = 12'h7D7;
        15'h0218: data = 12'h7DF;
        15'h0219: data = 12'h7E9;
        15'h021A: data = 12'h7EF;
        15'h021B: data = 12'h7F8;
        15'h021C: data = 12'h7FD;
        15'h021D: data = 12'h802;
        15'h021E: data = 12'h809;
        15'h021F: data = 12'h814;
        15'h0220: data = 12'h192;
        15'h0221: data = 12'h095;
        15'h0222: data = 12'h0A0;
        15'h0223: data = 12'h0A6;
        15'h0224: data = 12'h0A7;
        15'h0225: data = 12'h0B5;
        15'h0226: data = 12'h0B8;
        15'h0227: data = 12'h0BF;
        15'h0228: data = 12'h0BF;
        15'h0229: data = 12'h0C0;
        15'h022A: data = 12'h0C7;
        15'h022B: data = 12'h0C6;
        15'h022C: data = 12'h0C8;
        15'h022D: data = 12'h0C6;
        15'h022E: data = 12'h0CD;
        15'h022F: data = 12'h0CC;
        15'h0230: data = 12'h0C8;
        15'h0231: data = 12'h0C4;
        15'h0232: data = 12'h0C3;
        15'h0233: data = 12'h0C0;
        15'h0234: data = 12'h0C3;
        15'h0235: data = 12'h0BB;
        15'h0236: data = 12'h0BD;
        15'h0237: data = 12'h0C1;
        15'h0238: data = 12'h0C3;
        15'h0239: data = 12'h0C8;
        15'h023A: data = 12'h0C5;
        15'h023B: data = 12'h0C7;
        15'h023C: data = 12'h0C3;
        15'h023D: data = 12'h0C1;
        15'h023E: data = 12'h0B9;
        15'h023F: data = 12'h0B7;
        15'h0240: data = 12'h0AC;
        15'h0241: data = 12'h0A9;
        15'h0242: data = 12'h09D;
        15'h0243: data = 12'h095;
        15'h0244: data = 12'h094;
        15'h0245: data = 12'h091;
        15'h0246: data = 12'h08E;
        15'h0247: data = 12'h08D;
        15'h0248: data = 12'h088;
        15'h0249: data = 12'h086;
        15'h024A: data = 12'h07F;
        15'h024B: data = 12'h071;
        15'h024C: data = 12'h064;
        15'h024D: data = 12'h058;
        15'h024E: data = 12'h04C;
        15'h024F: data = 12'h04A;
        15'h0250: data = 12'h047;
        15'h0251: data = 12'h000;
        15'h0252: data = 12'h7C6;
        15'h0253: data = 12'h7BA;
        15'h0254: data = 12'h7AF;
        15'h0255: data = 12'h79F;
        15'h0256: data = 12'h789;
        15'h0257: data = 12'h77D;
        15'h0258: data = 12'h768;
        15'h0259: data = 12'h763;
        15'h025A: data = 12'h75D;
        15'h025B: data = 12'h758;
        15'h025C: data = 12'h74B;
        15'h025D: data = 12'h741;
        15'h025E: data = 12'h731;
        15'h025F: data = 12'h71F;
        15'h0260: data = 12'h70C;
        15'h0261: data = 12'h6FC;
        15'h0262: data = 12'h6ED;
        15'h0263: data = 12'h6DE;
        15'h0264: data = 12'h6DB;
        15'h0265: data = 12'h6CF;
        15'h0266: data = 12'h6C3;
        15'h0267: data = 12'h6B6;
        15'h0268: data = 12'h6A9;
        15'h0269: data = 12'h696;
        15'h026A: data = 12'h681;
        15'h026B: data = 12'h66B;
        15'h026C: data = 12'h657;
        15'h026D: data = 12'h647;
        15'h026E: data = 12'h637;
        15'h026F: data = 12'h62B;
        15'h0270: data = 12'h624;
        15'h0271: data = 12'h616;
        15'h0272: data = 12'h607;
        15'h0273: data = 12'h5F6;
        15'h0274: data = 12'h5DF;
        15'h0275: data = 12'h5D1;
        15'h0276: data = 12'h5C1;
        15'h0277: data = 12'h5B0;
        15'h0278: data = 12'h599;
        15'h0279: data = 12'h584;
        15'h027A: data = 12'h56A;
        15'h027B: data = 12'h556;
        15'h027C: data = 12'h543;
        15'h027D: data = 12'h52F;
        15'h027E: data = 12'h51C;
        15'h027F: data = 12'h50D;
        15'h0280: data = 12'h4FF;
        15'h0281: data = 12'h4E9;
        15'h0282: data = 12'h4D8;
        15'h0283: data = 12'h4CD;
        15'h0284: data = 12'h4B7;
        15'h0285: data = 12'h4A8;
        15'h0286: data = 12'h496;
        15'h0287: data = 12'h47C;
        15'h0288: data = 12'h466;
        15'h0289: data = 12'h456;
        15'h028A: data = 12'h440;
        15'h028B: data = 12'h427;
        15'h028C: data = 12'h40F;
        15'h028D: data = 12'h3F7;
        15'h028E: data = 12'h3E7;
        15'h028F: data = 12'h3D0;
        15'h0290: data = 12'h3B8;
        15'h0291: data = 12'h39C;
        15'h0292: data = 12'h388;
        15'h0293: data = 12'h36C;
        15'h0294: data = 12'h356;
        15'h0295: data = 12'h33B;
        15'h0296: data = 12'h32A;
        15'h0297: data = 12'h313;
        15'h0298: data = 12'h2FA;
        15'h0299: data = 12'h2E5;
        15'h029A: data = 12'h2CB;
        15'h029B: data = 12'h2B3;
        15'h029C: data = 12'h29C;
        15'h029D: data = 12'h283;
        15'h029E: data = 12'h26D;
        15'h029F: data = 12'h257;
        15'h02A0: data = 12'h23F;
        15'h02A1: data = 12'h22C;
        15'h02A2: data = 12'h20E;
        15'h02A3: data = 12'h1FC;
        15'h02A4: data = 12'h1E5;
        15'h02A5: data = 12'h1CB;
        15'h02A6: data = 12'h1AF;
        15'h02A7: data = 12'h19B;
        15'h02A8: data = 12'h183;
        15'h02A9: data = 12'h16D;
        15'h02AA: data = 12'h155;
        15'h02AB: data = 12'h140;
        15'h02AC: data = 12'h12A;
        15'h02AD: data = 12'h111;
        15'h02AE: data = 12'h0FA;
        15'h02AF: data = 12'h0E8;
        15'h02B0: data = 12'h0CE;
        15'h02B1: data = 12'h0B5;
        15'h02B2: data = 12'h097;
        15'h02B3: data = 12'h082;
        15'h02B4: data = 12'h075;
        15'h02B5: data = 12'h056;
        15'h02B6: data = 12'h03C;
        15'h02B7: data = 12'h7E2;
        15'h02B8: data = 12'h7C3;
        15'h02B9: data = 12'h7AA;
        15'h02BA: data = 12'h795;
        15'h02BB: data = 12'h780;
        15'h02BC: data = 12'h768;
        15'h02BD: data = 12'h751;
        15'h02BE: data = 12'h73E;
        15'h02BF: data = 12'h728;
        15'h02C0: data = 12'h711;
        15'h02C1: data = 12'h6F9;
        15'h02C2: data = 12'h6E4;
        15'h02C3: data = 12'h6D0;
        15'h02C4: data = 12'h6BC;
        15'h02C5: data = 12'h6A4;
        15'h02C6: data = 12'h68C;
        15'h02C7: data = 12'h680;
        15'h02C8: data = 12'h663;
        15'h02C9: data = 12'h655;
        15'h02CA: data = 12'h637;
        15'h02CB: data = 12'h628;
        15'h02CC: data = 12'h613;
        15'h02CD: data = 12'h5FF;
        15'h02CE: data = 12'h5E6;
        15'h02CF: data = 12'h5D0;
        15'h02D0: data = 12'h5C5;
        15'h02D1: data = 12'h5A9;
        15'h02D2: data = 12'h596;
        15'h02D3: data = 12'h57E;
        15'h02D4: data = 12'h56E;
        15'h02D5: data = 12'h55B;
        15'h02D6: data = 12'h544;
        15'h02D7: data = 12'h52C;
        15'h02D8: data = 12'h51F;
        15'h02D9: data = 12'h503;
        15'h02DA: data = 12'h4F0;
        15'h02DB: data = 12'h4E0;
        15'h02DC: data = 12'h4C7;
        15'h02DD: data = 12'h4B7;
        15'h02DE: data = 12'h4A0;
        15'h02DF: data = 12'h48B;
        15'h02E0: data = 12'h471;
        15'h02E1: data = 12'h45B;
        15'h02E2: data = 12'h447;
        15'h02E3: data = 12'h433;
        15'h02E4: data = 12'h41D;
        15'h02E5: data = 12'h40F;
        15'h02E6: data = 12'h3F5;
        15'h02E7: data = 12'h3E6;
        15'h02E8: data = 12'h3D8;
        15'h02E9: data = 12'h3C6;
        15'h02EA: data = 12'h3B3;
        15'h02EB: data = 12'h3A7;
        15'h02EC: data = 12'h399;
        15'h02ED: data = 12'h38D;
        15'h02EE: data = 12'h37E;
        15'h02EF: data = 12'h36D;
        15'h02F0: data = 12'h35E;
        15'h02F1: data = 12'h351;
        15'h02F2: data = 12'h342;
        15'h02F3: data = 12'h333;
        15'h02F4: data = 12'h322;
        15'h02F5: data = 12'h311;
        15'h02F6: data = 12'h2FE;
        15'h02F7: data = 12'h2EE;
        15'h02F8: data = 12'h2DB;
        15'h02F9: data = 12'h2CB;
        15'h02FA: data = 12'h2BA;
        15'h02FB: data = 12'h2AB;
        15'h02FC: data = 12'h299;
        15'h02FD: data = 12'h294;
        15'h02FE: data = 12'h285;
        15'h02FF: data = 12'h276;
        15'h0300: data = 12'h274;
        15'h0301: data = 12'h269;
        15'h0302: data = 12'h264;
        15'h0303: data = 12'h258;
        15'h0304: data = 12'h251;
        15'h0305: data = 12'h245;
        15'h0306: data = 12'h23B;
        15'h0307: data = 12'h228;
        15'h0308: data = 12'h21E;
        15'h0309: data = 12'h210;
        15'h030A: data = 12'h202;
        15'h030B: data = 12'h1F4;
        15'h030C: data = 12'h1E8;
        15'h030D: data = 12'h1E3;
        15'h030E: data = 12'h1DA;
        15'h030F: data = 12'h1D4;
        15'h0310: data = 12'h1D0;
        15'h0311: data = 12'h1C8;
        15'h0312: data = 12'h1C8;
        15'h0313: data = 12'h1C5;
        15'h0314: data = 12'h1BF;
        15'h0315: data = 12'h1B4;
        15'h0316: data = 12'h1AC;
        15'h0317: data = 12'h1A8;
        15'h0318: data = 12'h1A0;
        15'h0319: data = 12'h195;
        15'h031A: data = 12'h18A;
        15'h031B: data = 12'h187;
        15'h031C: data = 12'h17D;
        15'h031D: data = 12'h175;
        15'h031E: data = 12'h174;
        15'h031F: data = 12'h170;
        15'h0320: data = 12'h175;
        15'h0321: data = 12'h16F;
        15'h0322: data = 12'h175;
        15'h0323: data = 12'h179;
        15'h0324: data = 12'h16D;
        15'h0325: data = 12'h16F;
        15'h0326: data = 12'h16E;
        15'h0327: data = 12'h16D;
        15'h0328: data = 12'h163;
        15'h0329: data = 12'h15F;
        15'h032A: data = 12'h15D;
        15'h032B: data = 12'h157;
        15'h032C: data = 12'h155;
        15'h032D: data = 12'h154;
        15'h032E: data = 12'h156;
        15'h032F: data = 12'h15B;
        15'h0330: data = 12'h166;
        15'h0331: data = 12'h16A;
        15'h0332: data = 12'h16D;
        15'h0333: data = 12'h170;
        15'h0334: data = 12'h177;
        15'h0335: data = 12'h177;
        15'h0336: data = 12'h175;
        15'h0337: data = 12'h17E;
        15'h0338: data = 12'h17A;
        15'h0339: data = 12'h17F;
        15'h033A: data = 12'h17D;
        15'h033B: data = 12'h17D;
        15'h033C: data = 12'h185;
        15'h033D: data = 12'h181;
        15'h033E: data = 12'h18D;
        15'h033F: data = 12'h196;
        15'h0340: data = 12'h1A0;
        15'h0341: data = 12'h1AA;
        15'h0342: data = 12'h1B1;
        15'h0343: data = 12'h1BB;
        15'h0344: data = 12'h1C1;
        15'h0345: data = 12'h1CC;
        15'h0346: data = 12'h1D5;
        15'h0347: data = 12'h1DB;
        15'h0348: data = 12'h1E1;
        15'h0349: data = 12'h1E5;
        15'h034A: data = 12'h1E9;
        15'h034B: data = 12'h1ED;
        15'h034C: data = 12'h1F7;
        15'h034D: data = 12'h200;
        15'h034E: data = 12'h208;
        15'h034F: data = 12'h210;
        15'h0350: data = 12'h21F;
        15'h0351: data = 12'h226;
        15'h0352: data = 12'h239;
        15'h0353: data = 12'h247;
        15'h0354: data = 12'h25A;
        15'h0355: data = 12'h266;
        15'h0356: data = 12'h275;
        15'h0357: data = 12'h27D;
        15'h0358: data = 12'h28F;
        15'h0359: data = 12'h293;
        15'h035A: data = 12'h29F;
        15'h035B: data = 12'h2AF;
        15'h035C: data = 12'h2BB;
        15'h035D: data = 12'h2C2;
        15'h035E: data = 12'h2CD;
        15'h035F: data = 12'h2DB;
        15'h0360: data = 12'h2E6;
        15'h0361: data = 12'h2F7;
        15'h0362: data = 12'h305;
        15'h0363: data = 12'h317;
        15'h0364: data = 12'h329;
        15'h0365: data = 12'h339;
        15'h0366: data = 12'h34F;
        15'h0367: data = 12'h360;
        15'h0368: data = 12'h375;
        15'h0369: data = 12'h384;
        15'h036A: data = 12'h399;
        15'h036B: data = 12'h3A3;
        15'h036C: data = 12'h3BA;
        15'h036D: data = 12'h3C9;
        15'h036E: data = 12'h3D4;
        15'h036F: data = 12'h3EA;
        15'h0370: data = 12'h3F9;
        15'h0371: data = 12'h403;
        15'h0372: data = 12'h417;
        15'h0373: data = 12'h425;
        15'h0374: data = 12'h435;
        15'h0375: data = 12'h44A;
        15'h0376: data = 12'h45B;
        15'h0377: data = 12'h46F;
        15'h0378: data = 12'h482;
        15'h0379: data = 12'h49C;
        15'h037A: data = 12'h4AF;
        15'h037B: data = 12'h4C7;
        15'h037C: data = 12'h4DA;
        15'h037D: data = 12'h4F3;
        15'h037E: data = 12'h50B;
        15'h037F: data = 12'h51F;
        15'h0380: data = 12'h532;
        15'h0381: data = 12'h54B;
        15'h0382: data = 12'h561;
        15'h0383: data = 12'h573;
        15'h0384: data = 12'h581;
        15'h0385: data = 12'h595;
        15'h0386: data = 12'h5AA;
        15'h0387: data = 12'h5B8;
        15'h0388: data = 12'h5CD;
        15'h0389: data = 12'h5E2;
        15'h038A: data = 12'h5F5;
        15'h038B: data = 12'h60E;
        15'h038C: data = 12'h61C;
        15'h038D: data = 12'h634;
        15'h038E: data = 12'h651;
        15'h038F: data = 12'h663;
        15'h0390: data = 12'h683;
        15'h0391: data = 12'h698;
        15'h0392: data = 12'h6B3;
        15'h0393: data = 12'h6CC;
        15'h0394: data = 12'h6E4;
        15'h0395: data = 12'h6F9;
        15'h0396: data = 12'h714;
        15'h0397: data = 12'h72D;
        15'h0398: data = 12'h740;
        15'h0399: data = 12'h755;
        15'h039A: data = 12'h76E;
        15'h039B: data = 12'h784;
        15'h039C: data = 12'h79A;
        15'h039D: data = 12'h7AB;
        15'h039E: data = 12'h7C2;
        15'h039F: data = 12'h7D5;
        15'h03A0: data = 12'h7EA;
        15'h03A1: data = 12'h7FF;
        15'h03A2: data = 12'h064;
        15'h03A3: data = 12'h07D;
        15'h03A4: data = 12'h092;
        15'h03A5: data = 12'h0A4;
        15'h03A6: data = 12'h0BF;
        15'h03A7: data = 12'h0DB;
        15'h03A8: data = 12'h0F5;
        15'h03A9: data = 12'h107;
        15'h03AA: data = 12'h124;
        15'h03AB: data = 12'h140;
        15'h03AC: data = 12'h15A;
        15'h03AD: data = 12'h16C;
        15'h03AE: data = 12'h185;
        15'h03AF: data = 12'h1A0;
        15'h03B0: data = 12'h1BD;
        15'h03B1: data = 12'h1CB;
        15'h03B2: data = 12'h1E3;
        15'h03B3: data = 12'h1FB;
        15'h03B4: data = 12'h217;
        15'h03B5: data = 12'h224;
        15'h03B6: data = 12'h23D;
        15'h03B7: data = 12'h257;
        15'h03B8: data = 12'h26A;
        15'h03B9: data = 12'h279;
        15'h03BA: data = 12'h28D;
        15'h03BB: data = 12'h2A7;
        15'h03BC: data = 12'h2BD;
        15'h03BD: data = 12'h2CB;
        15'h03BE: data = 12'h2E9;
        15'h03BF: data = 12'h2FC;
        15'h03C0: data = 12'h318;
        15'h03C1: data = 12'h327;
        15'h03C2: data = 12'h33E;
        15'h03C3: data = 12'h356;
        15'h03C4: data = 12'h36C;
        15'h03C5: data = 12'h387;
        15'h03C6: data = 12'h39C;
        15'h03C7: data = 12'h3B4;
        15'h03C8: data = 12'h3D0;
        15'h03C9: data = 12'h3E3;
        15'h03CA: data = 12'h3F9;
        15'h03CB: data = 12'h410;
        15'h03CC: data = 12'h42D;
        15'h03CD: data = 12'h442;
        15'h03CE: data = 12'h453;
        15'h03CF: data = 12'h46A;
        15'h03D0: data = 12'h484;
        15'h03D1: data = 12'h497;
        15'h03D2: data = 12'h4AD;
        15'h03D3: data = 12'h4BF;
        15'h03D4: data = 12'h4D4;
        15'h03D5: data = 12'h4E8;
        15'h03D6: data = 12'h4FD;
        15'h03D7: data = 12'h511;
        15'h03D8: data = 12'h51B;
        15'h03D9: data = 12'h534;
        15'h03DA: data = 12'h54B;
        15'h03DB: data = 12'h556;
        15'h03DC: data = 12'h56D;
        15'h03DD: data = 12'h579;
        15'h03DE: data = 12'h58E;
        15'h03DF: data = 12'h5A0;
        15'h03E0: data = 12'h5AF;
        15'h03E1: data = 12'h5C4;
        15'h03E2: data = 12'h5CD;
        15'h03E3: data = 12'h5DE;
        15'h03E4: data = 12'h5EE;
        15'h03E5: data = 12'h5FF;
        15'h03E6: data = 12'h611;
        15'h03E7: data = 12'h61A;
        15'h03E8: data = 12'h62B;
        15'h03E9: data = 12'h638;
        15'h03EA: data = 12'h648;
        15'h03EB: data = 12'h65E;
        15'h03EC: data = 12'h66C;
        15'h03ED: data = 12'h675;
        15'h03EE: data = 12'h688;
        15'h03EF: data = 12'h697;
        15'h03F0: data = 12'h6A4;
        15'h03F1: data = 12'h6B7;
        15'h03F2: data = 12'h6C1;
        15'h03F3: data = 12'h6CC;
        15'h03F4: data = 12'h6E1;
        15'h03F5: data = 12'h6EE;
        15'h03F6: data = 12'h6F2;
        15'h03F7: data = 12'h708;
        15'h03F8: data = 12'h718;
        15'h03F9: data = 12'h725;
        15'h03FA: data = 12'h72E;
        15'h03FB: data = 12'h735;
        15'h03FC: data = 12'h741;
        15'h03FD: data = 12'h756;
        15'h03FE: data = 12'h75F;
        15'h03FF: data = 12'h76D;
        15'h0400: data = 12'h778;
        15'h0401: data = 12'h785;
        15'h0402: data = 12'h790;
        15'h0403: data = 12'h79A;
        15'h0404: data = 12'h7A4;
        15'h0405: data = 12'h7AF;
        15'h0406: data = 12'h7B8;
        15'h0407: data = 12'h7BF;
        15'h0408: data = 12'h7C8;
        15'h0409: data = 12'h7CF;
        15'h040A: data = 12'h7DA;
        15'h040B: data = 12'h7E0;
        15'h040C: data = 12'h7EA;
        15'h040D: data = 12'h7F2;
        15'h040E: data = 12'h7F7;
        15'h040F: data = 12'h7FD;
        15'h0410: data = 12'h807;
        15'h0411: data = 12'h807;
        15'h0412: data = 12'h80E;
        15'h0413: data = 12'h818;
        15'h0414: data = 12'h096;
        15'h0415: data = 12'h09A;
        15'h0416: data = 12'h0A2;
        15'h0417: data = 12'h0A5;
        15'h0418: data = 12'h0A8;
        15'h0419: data = 12'h0B0;
        15'h041A: data = 12'h0B2;
        15'h041B: data = 12'h0BC;
        15'h041C: data = 12'h0BA;
        15'h041D: data = 12'h0B9;
        15'h041E: data = 12'h0BC;
        15'h041F: data = 12'h0BE;
        15'h0420: data = 12'h0BB;
        15'h0421: data = 12'h0B8;
        15'h0422: data = 12'h0C1;
        15'h0423: data = 12'h0C1;
        15'h0424: data = 12'h0C5;
        15'h0425: data = 12'h0C3;
        15'h0426: data = 12'h0C6;
        15'h0427: data = 12'h0C8;
        15'h0428: data = 12'h0CD;
        15'h0429: data = 12'h0C8;
        15'h042A: data = 12'h0CC;
        15'h042B: data = 12'h0D0;
        15'h042C: data = 12'h0CF;
        15'h042D: data = 12'h0D0;
        15'h042E: data = 12'h0C8;
        15'h042F: data = 12'h0C9;
        15'h0430: data = 12'h0BD;
        15'h0431: data = 12'h0B8;
        15'h0432: data = 12'h0AE;
        15'h0433: data = 12'h0A8;
        15'h0434: data = 12'h0A3;
        15'h0435: data = 12'h0A4;
        15'h0436: data = 12'h0A0;
        15'h0437: data = 12'h09F;
        15'h0438: data = 12'h0A4;
        15'h0439: data = 12'h09F;
        15'h043A: data = 12'h098;
        15'h043B: data = 12'h091;
        15'h043C: data = 12'h086;
        15'h043D: data = 12'h07D;
        15'h043E: data = 12'h072;
        15'h043F: data = 12'h069;
        15'h0440: data = 12'h061;
        15'h0441: data = 12'h05C;
        15'h0442: data = 12'h05E;
        15'h0443: data = 12'h05A;
        15'h0444: data = 12'h054;
        15'h0445: data = 12'h042;
        15'h0446: data = 12'h7C2;
        15'h0447: data = 12'h7B1;
        15'h0448: data = 12'h7A2;
        15'h0449: data = 12'h795;
        15'h044A: data = 12'h784;
        15'h044B: data = 12'h785;
        15'h044C: data = 12'h77B;
        15'h044D: data = 12'h775;
        15'h044E: data = 12'h765;
        15'h044F: data = 12'h756;
        15'h0450: data = 12'h744;
        15'h0451: data = 12'h732;
        15'h0452: data = 12'h722;
        15'h0453: data = 12'h719;
        15'h0454: data = 12'h70C;
        15'h0455: data = 12'h704;
        15'h0456: data = 12'h6F9;
        15'h0457: data = 12'h6EC;
        15'h0458: data = 12'h6E4;
        15'h0459: data = 12'h6D5;
        15'h045A: data = 12'h6BF;
        15'h045B: data = 12'h6AF;
        15'h045C: data = 12'h699;
        15'h045D: data = 12'h685;
        15'h045E: data = 12'h678;
        15'h045F: data = 12'h66B;
        15'h0460: data = 12'h65D;
        15'h0461: data = 12'h656;
        15'h0462: data = 12'h64A;
        15'h0463: data = 12'h63B;
        15'h0464: data = 12'h62F;
        15'h0465: data = 12'h617;
        15'h0466: data = 12'h605;
        15'h0467: data = 12'h5F2;
        15'h0468: data = 12'h5D7;
        15'h0469: data = 12'h5C3;
        15'h046A: data = 12'h5B3;
        15'h046B: data = 12'h5A2;
        15'h046C: data = 12'h58E;
        15'h046D: data = 12'h57D;
        15'h046E: data = 12'h568;
        15'h046F: data = 12'h55D;
        15'h0470: data = 12'h552;
        15'h0471: data = 12'h540;
        15'h0472: data = 12'h52C;
        15'h0473: data = 12'h521;
        15'h0474: data = 12'h50E;
        15'h0475: data = 12'h4F5;
        15'h0476: data = 12'h4DD;
        15'h0477: data = 12'h4CE;
        15'h0478: data = 12'h4B8;
        15'h0479: data = 12'h49F;
        15'h047A: data = 12'h488;
        15'h047B: data = 12'h471;
        15'h047C: data = 12'h45B;
        15'h047D: data = 12'h448;
        15'h047E: data = 12'h42E;
        15'h047F: data = 12'h417;
        15'h0480: data = 12'h3FF;
        15'h0481: data = 12'h3E5;
        15'h0482: data = 12'h3D7;
        15'h0483: data = 12'h3C3;
        15'h0484: data = 12'h3AD;
        15'h0485: data = 12'h395;
        15'h0486: data = 12'h383;
        15'h0487: data = 12'h368;
        15'h0488: data = 12'h357;
        15'h0489: data = 12'h33D;
        15'h048A: data = 12'h32D;
        15'h048B: data = 12'h319;
        15'h048C: data = 12'h301;
        15'h048D: data = 12'h2EE;
        15'h048E: data = 12'h2D5;
        15'h048F: data = 12'h2C1;
        15'h0490: data = 12'h2AC;
        15'h0491: data = 12'h291;
        15'h0492: data = 12'h27C;
        15'h0493: data = 12'h267;
        15'h0494: data = 12'h24E;
        15'h0495: data = 12'h23A;
        15'h0496: data = 12'h21D;
        15'h0497: data = 12'h20A;
        15'h0498: data = 12'h1F5;
        15'h0499: data = 12'h1DD;
        15'h049A: data = 12'h1C1;
        15'h049B: data = 12'h1AB;
        15'h049C: data = 12'h197;
        15'h049D: data = 12'h17E;
        15'h049E: data = 12'h165;
        15'h049F: data = 12'h14F;
        15'h04A0: data = 12'h138;
        15'h04A1: data = 12'h11E;
        15'h04A2: data = 12'h109;
        15'h04A3: data = 12'h0F6;
        15'h04A4: data = 12'h0DD;
        15'h04A5: data = 12'h0C3;
        15'h04A6: data = 12'h0AB;
        15'h04A7: data = 12'h093;
        15'h04A8: data = 12'h085;
        15'h04A9: data = 12'h06A;
        15'h04AA: data = 12'h04E;
        15'h04AB: data = 12'h3A1;
        15'h04AC: data = 12'h7D4;
        15'h04AD: data = 12'h7BB;
        15'h04AE: data = 12'h7A2;
        15'h04AF: data = 12'h78C;
        15'h04B0: data = 12'h778;
        15'h04B1: data = 12'h762;
        15'h04B2: data = 12'h74C;
        15'h04B3: data = 12'h739;
        15'h04B4: data = 12'h71C;
        15'h04B5: data = 12'h708;
        15'h04B6: data = 12'h6F3;
        15'h04B7: data = 12'h6DC;
        15'h04B8: data = 12'h6CA;
        15'h04B9: data = 12'h6B1;
        15'h04BA: data = 12'h699;
        15'h04BB: data = 12'h68A;
        15'h04BC: data = 12'h66C;
        15'h04BD: data = 12'h65C;
        15'h04BE: data = 12'h640;
        15'h04BF: data = 12'h630;
        15'h04C0: data = 12'h617;
        15'h04C1: data = 12'h5FE;
        15'h04C2: data = 12'h5EA;
        15'h04C3: data = 12'h5CF;
        15'h04C4: data = 12'h5BF;
        15'h04C5: data = 12'h5A4;
        15'h04C6: data = 12'h591;
        15'h04C7: data = 12'h579;
        15'h04C8: data = 12'h56A;
        15'h04C9: data = 12'h556;
        15'h04CA: data = 12'h539;
        15'h04CB: data = 12'h524;
        15'h04CC: data = 12'h513;
        15'h04CD: data = 12'h4F9;
        15'h04CE: data = 12'h4E3;
        15'h04CF: data = 12'h4D0;
        15'h04D0: data = 12'h4B6;
        15'h04D1: data = 12'h4A7;
        15'h04D2: data = 12'h492;
        15'h04D3: data = 12'h481;
        15'h04D4: data = 12'h467;
        15'h04D5: data = 12'h455;
        15'h04D6: data = 12'h446;
        15'h04D7: data = 12'h438;
        15'h04D8: data = 12'h420;
        15'h04D9: data = 12'h417;
        15'h04DA: data = 12'h3FF;
        15'h04DB: data = 12'h3F6;
        15'h04DC: data = 12'h3E7;
        15'h04DD: data = 12'h3D5;
        15'h04DE: data = 12'h3C6;
        15'h04DF: data = 12'h3B7;
        15'h04E0: data = 12'h3A5;
        15'h04E1: data = 12'h396;
        15'h04E2: data = 12'h37E;
        15'h04E3: data = 12'h36B;
        15'h04E4: data = 12'h35A;
        15'h04E5: data = 12'h344;
        15'h04E6: data = 12'h336;
        15'h04E7: data = 12'h327;
        15'h04E8: data = 12'h314;
        15'h04E9: data = 12'h300;
        15'h04EA: data = 12'h2EF;
        15'h04EB: data = 12'h2E1;
        15'h04EC: data = 12'h2D5;
        15'h04ED: data = 12'h2CD;
        15'h04EE: data = 12'h2BF;
        15'h04EF: data = 12'h2B7;
        15'h04F0: data = 12'h2A9;
        15'h04F1: data = 12'h2A0;
        15'h04F2: data = 12'h296;
        15'h04F3: data = 12'h283;
        15'h04F4: data = 12'h27F;
        15'h04F5: data = 12'h26D;
        15'h04F6: data = 12'h265;
        15'h04F7: data = 12'h251;
        15'h04F8: data = 12'h249;
        15'h04F9: data = 12'h232;
        15'h04FA: data = 12'h229;
        15'h04FB: data = 12'h219;
        15'h04FC: data = 12'h210;
        15'h04FD: data = 12'h207;
        15'h04FE: data = 12'h200;
        15'h04FF: data = 12'h1F4;
        15'h0500: data = 12'h1EF;
        15'h0501: data = 12'h1EC;
        15'h0502: data = 12'h1E8;
        15'h0503: data = 12'h1E2;
        15'h0504: data = 12'h1DF;
        15'h0505: data = 12'h1D0;
        15'h0506: data = 12'h1CA;
        15'h0507: data = 12'h1C3;
        15'h0508: data = 12'h1B5;
        15'h0509: data = 12'h1AB;
        15'h050A: data = 12'h19F;
        15'h050B: data = 12'h197;
        15'h050C: data = 12'h191;
        15'h050D: data = 12'h18A;
        15'h050E: data = 12'h183;
        15'h050F: data = 12'h188;
        15'h0510: data = 12'h186;
        15'h0511: data = 12'h182;
        15'h0512: data = 12'h183;
        15'h0513: data = 12'h17C;
        15'h0514: data = 12'h181;
        15'h0515: data = 12'h176;
        15'h0516: data = 12'h176;
        15'h0517: data = 12'h175;
        15'h0518: data = 12'h167;
        15'h0519: data = 12'h166;
        15'h051A: data = 12'h162;
        15'h051B: data = 12'h15C;
        15'h051C: data = 12'h157;
        15'h051D: data = 12'h152;
        15'h051E: data = 12'h157;
        15'h051F: data = 12'h15A;
        15'h0520: data = 12'h15E;
        15'h0521: data = 12'h163;
        15'h0522: data = 12'h165;
        15'h0523: data = 12'h16B;
        15'h0524: data = 12'h16F;
        15'h0525: data = 12'h16C;
        15'h0526: data = 12'h16E;
        15'h0527: data = 12'h16B;
        15'h0528: data = 12'h16F;
        15'h0529: data = 12'h16C;
        15'h052A: data = 12'h167;
        15'h052B: data = 12'h16E;
        15'h052C: data = 12'h16A;
        15'h052D: data = 12'h176;
        15'h052E: data = 12'h177;
        15'h052F: data = 12'h17E;
        15'h0530: data = 12'h18E;
        15'h0531: data = 12'h18E;
        15'h0532: data = 12'h19C;
        15'h0533: data = 12'h1A6;
        15'h0534: data = 12'h1A9;
        15'h0535: data = 12'h1AF;
        15'h0536: data = 12'h1B1;
        15'h0537: data = 12'h1BA;
        15'h0538: data = 12'h1C1;
        15'h0539: data = 12'h1C2;
        15'h053A: data = 12'h1C5;
        15'h053B: data = 12'h1CA;
        15'h053C: data = 12'h1CD;
        15'h053D: data = 12'h1D6;
        15'h053E: data = 12'h1DF;
        15'h053F: data = 12'h1E9;
        15'h0540: data = 12'h1F9;
        15'h0541: data = 12'h206;
        15'h0542: data = 12'h213;
        15'h0543: data = 12'h21C;
        15'h0544: data = 12'h230;
        15'h0545: data = 12'h238;
        15'h0546: data = 12'h242;
        15'h0547: data = 12'h24D;
        15'h0548: data = 12'h25B;
        15'h0549: data = 12'h261;
        15'h054A: data = 12'h26F;
        15'h054B: data = 12'h273;
        15'h054C: data = 12'h282;
        15'h054D: data = 12'h285;
        15'h054E: data = 12'h291;
        15'h054F: data = 12'h2A3;
        15'h0550: data = 12'h2AE;
        15'h0551: data = 12'h2BE;
        15'h0552: data = 12'h2C9;
        15'h0553: data = 12'h2DE;
        15'h0554: data = 12'h2F0;
        15'h0555: data = 12'h303;
        15'h0556: data = 12'h318;
        15'h0557: data = 12'h326;
        15'h0558: data = 12'h336;
        15'h0559: data = 12'h344;
        15'h055A: data = 12'h356;
        15'h055B: data = 12'h365;
        15'h055C: data = 12'h372;
        15'h055D: data = 12'h380;
        15'h055E: data = 12'h394;
        15'h055F: data = 12'h397;
        15'h0560: data = 12'h3A8;
        15'h0561: data = 12'h3B9;
        15'h0562: data = 12'h3C6;
        15'h0563: data = 12'h3D8;
        15'h0564: data = 12'h3EC;
        15'h0565: data = 12'h3FE;
        15'h0566: data = 12'h414;
        15'h0567: data = 12'h428;
        15'h0568: data = 12'h43D;
        15'h0569: data = 12'h454;
        15'h056A: data = 12'h469;
        15'h056B: data = 12'h480;
        15'h056C: data = 12'h490;
        15'h056D: data = 12'h4AA;
        15'h056E: data = 12'h4B8;
        15'h056F: data = 12'h4CF;
        15'h0570: data = 12'h4DC;
        15'h0571: data = 12'h4F1;
        15'h0572: data = 12'h505;
        15'h0573: data = 12'h517;
        15'h0574: data = 12'h52E;
        15'h0575: data = 12'h53D;
        15'h0576: data = 12'h553;
        15'h0577: data = 12'h561;
        15'h0578: data = 12'h572;
        15'h0579: data = 12'h586;
        15'h057A: data = 12'h599;
        15'h057B: data = 12'h5B4;
        15'h057C: data = 12'h5CA;
        15'h057D: data = 12'h5E5;
        15'h057E: data = 12'h600;
        15'h057F: data = 12'h618;
        15'h0580: data = 12'h62D;
        15'h0581: data = 12'h646;
        15'h0582: data = 12'h65F;
        15'h0583: data = 12'h676;
        15'h0584: data = 12'h690;
        15'h0585: data = 12'h6A0;
        15'h0586: data = 12'h6B8;
        15'h0587: data = 12'h6CF;
        15'h0588: data = 12'h6E1;
        15'h0589: data = 12'h6F4;
        15'h058A: data = 12'h70C;
        15'h058B: data = 12'h720;
        15'h058C: data = 12'h732;
        15'h058D: data = 12'h746;
        15'h058E: data = 12'h75D;
        15'h058F: data = 12'h773;
        15'h0590: data = 12'h788;
        15'h0591: data = 12'h79E;
        15'h0592: data = 12'h7B7;
        15'h0593: data = 12'h7CE;
        15'h0594: data = 12'h7E4;
        15'h0595: data = 12'h7FF;
        15'h0596: data = 12'h136;
        15'h0597: data = 12'h087;
        15'h0598: data = 12'h09D;
        15'h0599: data = 12'h0B0;
        15'h059A: data = 12'h0CD;
        15'h059B: data = 12'h0E6;
        15'h059C: data = 12'h100;
        15'h059D: data = 12'h111;
        15'h059E: data = 12'h12C;
        15'h059F: data = 12'h144;
        15'h05A0: data = 12'h155;
        15'h05A1: data = 12'h16B;
        15'h05A2: data = 12'h17F;
        15'h05A3: data = 12'h197;
        15'h05A4: data = 12'h1B0;
        15'h05A5: data = 12'h1C0;
        15'h05A6: data = 12'h1D7;
        15'h05A7: data = 12'h1EF;
        15'h05A8: data = 12'h207;
        15'h05A9: data = 12'h218;
        15'h05AA: data = 12'h230;
        15'h05AB: data = 12'h24A;
        15'h05AC: data = 12'h261;
        15'h05AD: data = 12'h274;
        15'h05AE: data = 12'h287;
        15'h05AF: data = 12'h2A6;
        15'h05B0: data = 12'h2C1;
        15'h05B1: data = 12'h2D5;
        15'h05B2: data = 12'h2F2;
        15'h05B3: data = 12'h308;
        15'h05B4: data = 12'h325;
        15'h05B5: data = 12'h334;
        15'h05B6: data = 12'h34F;
        15'h05B7: data = 12'h366;
        15'h05B8: data = 12'h37B;
        15'h05B9: data = 12'h395;
        15'h05BA: data = 12'h3A8;
        15'h05BB: data = 12'h3C1;
        15'h05BC: data = 12'h3DB;
        15'h05BD: data = 12'h3F0;
        15'h05BE: data = 12'h3FF;
        15'h05BF: data = 12'h417;
        15'h05C0: data = 12'h42F;
        15'h05C1: data = 12'h443;
        15'h05C2: data = 12'h454;
        15'h05C3: data = 12'h469;
        15'h05C4: data = 12'h480;
        15'h05C5: data = 12'h493;
        15'h05C6: data = 12'h4A6;
        15'h05C7: data = 12'h4B8;
        15'h05C8: data = 12'h4C9;
        15'h05C9: data = 12'h4DB;
        15'h05CA: data = 12'h4F1;
        15'h05CB: data = 12'h503;
        15'h05CC: data = 12'h50E;
        15'h05CD: data = 12'h525;
        15'h05CE: data = 12'h53D;
        15'h05CF: data = 12'h546;
        15'h05D0: data = 12'h55B;
        15'h05D1: data = 12'h56A;
        15'h05D2: data = 12'h580;
        15'h05D3: data = 12'h590;
        15'h05D4: data = 12'h5A3;
        15'h05D5: data = 12'h5B6;
        15'h05D6: data = 12'h5C6;
        15'h05D7: data = 12'h5D4;
        15'h05D8: data = 12'h5E8;
        15'h05D9: data = 12'h5FD;
        15'h05DA: data = 12'h60C;
        15'h05DB: data = 12'h61D;
        15'h05DC: data = 12'h62D;
        15'h05DD: data = 12'h63B;
        15'h05DE: data = 12'h64F;
        15'h05DF: data = 12'h660;
        15'h05E0: data = 12'h671;
        15'h05E1: data = 12'h67F;
        15'h05E2: data = 12'h695;
        15'h05E3: data = 12'h6A1;
        15'h05E4: data = 12'h6AF;
        15'h05E5: data = 12'h6C2;
        15'h05E6: data = 12'h6D1;
        15'h05E7: data = 12'h6DC;
        15'h05E8: data = 12'h6EC;
        15'h05E9: data = 12'h6FA;
        15'h05EA: data = 12'h705;
        15'h05EB: data = 12'h716;
        15'h05EC: data = 12'h725;
        15'h05ED: data = 12'h732;
        15'h05EE: data = 12'h738;
        15'h05EF: data = 12'h744;
        15'h05F0: data = 12'h752;
        15'h05F1: data = 12'h761;
        15'h05F2: data = 12'h768;
        15'h05F3: data = 12'h779;
        15'h05F4: data = 12'h77F;
        15'h05F5: data = 12'h78D;
        15'h05F6: data = 12'h799;
        15'h05F7: data = 12'h79B;
        15'h05F8: data = 12'h7A2;
        15'h05F9: data = 12'h7AD;
        15'h05FA: data = 12'h7B8;
        15'h05FB: data = 12'h7C0;
        15'h05FC: data = 12'h7C9;
        15'h05FD: data = 12'h7CD;
        15'h05FE: data = 12'h7D2;
        15'h05FF: data = 12'h7DC;
        15'h0600: data = 12'h7E3;
        15'h0601: data = 12'h7EB;
        15'h0602: data = 12'h7F2;
        15'h0603: data = 12'h7F6;
        15'h0604: data = 12'h7FF;
        15'h0605: data = 12'h7FF;
        15'h0606: data = 12'h802;
        15'h0607: data = 12'h80D;
        15'h0608: data = 12'h7ED;
        15'h0609: data = 12'h089;
        15'h060A: data = 12'h092;
        15'h060B: data = 12'h097;
        15'h060C: data = 12'h098;
        15'h060D: data = 12'h0A0;
        15'h060E: data = 12'h0A4;
        15'h060F: data = 12'h0AD;
        15'h0610: data = 12'h0AD;
        15'h0611: data = 12'h0AD;
        15'h0612: data = 12'h0B5;
        15'h0613: data = 12'h0B7;
        15'h0614: data = 12'h0BA;
        15'h0615: data = 12'h0B9;
        15'h0616: data = 12'h0C3;
        15'h0617: data = 12'h0C7;
        15'h0618: data = 12'h0CC;
        15'h0619: data = 12'h0D0;
        15'h061A: data = 12'h0D1;
        15'h061B: data = 12'h0D5;
        15'h061C: data = 12'h0D6;
        15'h061D: data = 12'h0CD;
        15'h061E: data = 12'h0CF;
        15'h061F: data = 12'h0CB;
        15'h0620: data = 12'h0CC;
        15'h0621: data = 12'h0C7;
        15'h0622: data = 12'h0BC;
        15'h0623: data = 12'h0B6;
        15'h0624: data = 12'h0AF;
        15'h0625: data = 12'h0AF;
        15'h0626: data = 12'h0A6;
        15'h0627: data = 12'h0A9;
        15'h0628: data = 12'h0AA;
        15'h0629: data = 12'h0B1;
        15'h062A: data = 12'h0AB;
        15'h062B: data = 12'h0A7;
        15'h062C: data = 12'h0A6;
        15'h062D: data = 12'h09A;
        15'h062E: data = 12'h090;
        15'h062F: data = 12'h081;
        15'h0630: data = 12'h077;
        15'h0631: data = 12'h078;
        15'h0632: data = 12'h06D;
        15'h0633: data = 12'h06A;
        15'h0634: data = 12'h069;
        15'h0635: data = 12'h068;
        15'h0636: data = 12'h061;
        15'h0637: data = 12'h059;
        15'h0638: data = 12'h04D;
        15'h0639: data = 12'h038;
        15'h063A: data = 12'h7B5;
        15'h063B: data = 12'h7A8;
        15'h063C: data = 12'h7A3;
        15'h063D: data = 12'h79C;
        15'h063E: data = 12'h794;
        15'h063F: data = 12'h78D;
        15'h0640: data = 12'h77F;
        15'h0641: data = 12'h772;
        15'h0642: data = 12'h75E;
        15'h0643: data = 12'h74B;
        15'h0644: data = 12'h739;
        15'h0645: data = 12'h731;
        15'h0646: data = 12'h724;
        15'h0647: data = 12'h71E;
        15'h0648: data = 12'h71B;
        15'h0649: data = 12'h70D;
        15'h064A: data = 12'h6FC;
        15'h064B: data = 12'h6EA;
        15'h064C: data = 12'h6DE;
        15'h064D: data = 12'h6CB;
        15'h064E: data = 12'h6B3;
        15'h064F: data = 12'h6A3;
        15'h0650: data = 12'h694;
        15'h0651: data = 12'h689;
        15'h0652: data = 12'h67D;
        15'h0653: data = 12'h676;
        15'h0654: data = 12'h666;
        15'h0655: data = 12'h65A;
        15'h0656: data = 12'h647;
        15'h0657: data = 12'h634;
        15'h0658: data = 12'h62A;
        15'h0659: data = 12'h60E;
        15'h065A: data = 12'h5F7;
        15'h065B: data = 12'h5E3;
        15'h065C: data = 12'h5D0;
        15'h065D: data = 12'h5BB;
        15'h065E: data = 12'h5B2;
        15'h065F: data = 12'h5A5;
        15'h0660: data = 12'h594;
        15'h0661: data = 12'h586;
        15'h0662: data = 12'h571;
        15'h0663: data = 12'h564;
        15'h0664: data = 12'h559;
        15'h0665: data = 12'h544;
        15'h0666: data = 12'h52B;
        15'h0667: data = 12'h51B;
        15'h0668: data = 12'h50A;
        15'h0669: data = 12'h4F6;
        15'h066A: data = 12'h4D5;
        15'h066B: data = 12'h4C5;
        15'h066C: data = 12'h4AB;
        15'h066D: data = 12'h498;
        15'h066E: data = 12'h47F;
        15'h066F: data = 12'h467;
        15'h0670: data = 12'h454;
        15'h0671: data = 12'h445;
        15'h0672: data = 12'h42F;
        15'h0673: data = 12'h417;
        15'h0674: data = 12'h3FF;
        15'h0675: data = 12'h3EB;
        15'h0676: data = 12'h3DA;
        15'h0677: data = 12'h3C6;
        15'h0678: data = 12'h3B1;
        15'h0679: data = 12'h39C;
        15'h067A: data = 12'h38B;
        15'h067B: data = 12'h370;
        15'h067C: data = 12'h35D;
        15'h067D: data = 12'h344;
        15'h067E: data = 12'h338;
        15'h067F: data = 12'h322;
        15'h0680: data = 12'h306;
        15'h0681: data = 12'h2F4;
        15'h0682: data = 12'h2DD;
        15'h0683: data = 12'h2C7;
        15'h0684: data = 12'h2AE;
        15'h0685: data = 12'h295;
        15'h0686: data = 12'h27E;
        15'h0687: data = 12'h26D;
        15'h0688: data = 12'h250;
        15'h0689: data = 12'h23E;
        15'h068A: data = 12'h221;
        15'h068B: data = 12'h20D;
        15'h068C: data = 12'h1F6;
        15'h068D: data = 12'h1DC;
        15'h068E: data = 12'h1C4;
        15'h068F: data = 12'h1AC;
        15'h0690: data = 12'h199;
        15'h0691: data = 12'h17F;
        15'h0692: data = 12'h167;
        15'h0693: data = 12'h14D;
        15'h0694: data = 12'h13B;
        15'h0695: data = 12'h11E;
        15'h0696: data = 12'h108;
        15'h0697: data = 12'h0F4;
        15'h0698: data = 12'h0DD;
        15'h0699: data = 12'h0C4;
        15'h069A: data = 12'h0AA;
        15'h069B: data = 12'h098;
        15'h069C: data = 12'h084;
        15'h069D: data = 12'h066;
        15'h069E: data = 12'h04C;
        15'h069F: data = 12'h7E0;
        15'h06A0: data = 12'h7D1;
        15'h06A1: data = 12'h7B9;
        15'h06A2: data = 12'h7A2;
        15'h06A3: data = 12'h78C;
        15'h06A4: data = 12'h775;
        15'h06A5: data = 12'h75F;
        15'h06A6: data = 12'h74A;
        15'h06A7: data = 12'h732;
        15'h06A8: data = 12'h71A;
        15'h06A9: data = 12'h704;
        15'h06AA: data = 12'h6ED;
        15'h06AB: data = 12'h6D5;
        15'h06AC: data = 12'h6C0;
        15'h06AD: data = 12'h6A9;
        15'h06AE: data = 12'h694;
        15'h06AF: data = 12'h684;
        15'h06B0: data = 12'h669;
        15'h06B1: data = 12'h654;
        15'h06B2: data = 12'h639;
        15'h06B3: data = 12'h626;
        15'h06B4: data = 12'h612;
        15'h06B5: data = 12'h5F7;
        15'h06B6: data = 12'h5E0;
        15'h06B7: data = 12'h5C6;
        15'h06B8: data = 12'h5B8;
        15'h06B9: data = 12'h59A;
        15'h06BA: data = 12'h584;
        15'h06BB: data = 12'h56B;
        15'h06BC: data = 12'h55D;
        15'h06BD: data = 12'h549;
        15'h06BE: data = 12'h531;
        15'h06BF: data = 12'h51D;
        15'h06C0: data = 12'h50B;
        15'h06C1: data = 12'h4F2;
        15'h06C2: data = 12'h4E0;
        15'h06C3: data = 12'h4CF;
        15'h06C4: data = 12'h4B7;
        15'h06C5: data = 12'h4A8;
        15'h06C6: data = 12'h493;
        15'h06C7: data = 12'h487;
        15'h06C8: data = 12'h471;
        15'h06C9: data = 12'h460;
        15'h06CA: data = 12'h450;
        15'h06CB: data = 12'h441;
        15'h06CC: data = 12'h42C;
        15'h06CD: data = 12'h420;
        15'h06CE: data = 12'h407;
        15'h06CF: data = 12'h3FB;
        15'h06D0: data = 12'h3E9;
        15'h06D1: data = 12'h3D3;
        15'h06D2: data = 12'h3BD;
        15'h06D3: data = 12'h3B0;
        15'h06D4: data = 12'h39B;
        15'h06D5: data = 12'h38E;
        15'h06D6: data = 12'h376;
        15'h06D7: data = 12'h362;
        15'h06D8: data = 12'h34E;
        15'h06D9: data = 12'h33E;
        15'h06DA: data = 12'h32F;
        15'h06DB: data = 12'h31F;
        15'h06DC: data = 12'h30F;
        15'h06DD: data = 12'h300;
        15'h06DE: data = 12'h2F4;
        15'h06DF: data = 12'h2E8;
        15'h06E0: data = 12'h2DD;
        15'h06E1: data = 12'h2DA;
        15'h06E2: data = 12'h2C8;
        15'h06E3: data = 12'h2BB;
        15'h06E4: data = 12'h2AF;
        15'h06E5: data = 12'h2A1;
        15'h06E6: data = 12'h295;
        15'h06E7: data = 12'h284;
        15'h06E8: data = 12'h277;
        15'h06E9: data = 12'h267;
        15'h06EA: data = 12'h25B;
        15'h06EB: data = 12'h247;
        15'h06EC: data = 12'h23E;
        15'h06ED: data = 12'h22D;
        15'h06EE: data = 12'h227;
        15'h06EF: data = 12'h216;
        15'h06F0: data = 12'h212;
        15'h06F1: data = 12'h20E;
        15'h06F2: data = 12'h20A;
        15'h06F3: data = 12'h200;
        15'h06F4: data = 12'h1F7;
        15'h06F5: data = 12'h1F3;
        15'h06F6: data = 12'h1ED;
        15'h06F7: data = 12'h1E4;
        15'h06F8: data = 12'h1D7;
        15'h06F9: data = 12'h1C9;
        15'h06FA: data = 12'h1C1;
        15'h06FB: data = 12'h1B6;
        15'h06FC: data = 12'h1AB;
        15'h06FD: data = 12'h1A0;
        15'h06FE: data = 12'h19C;
        15'h06FF: data = 12'h199;
        15'h0700: data = 12'h196;
        15'h0701: data = 12'h193;
        15'h0702: data = 12'h191;
        15'h0703: data = 12'h192;
        15'h0704: data = 12'h18F;
        15'h0705: data = 12'h189;
        15'h0706: data = 12'h185;
        15'h0707: data = 12'h180;
        15'h0708: data = 12'h17A;
        15'h0709: data = 12'h175;
        15'h070A: data = 12'h16F;
        15'h070B: data = 12'h16A;
        15'h070C: data = 12'h161;
        15'h070D: data = 12'h15E;
        15'h070E: data = 12'h15C;
        15'h070F: data = 12'h15F;
        15'h0710: data = 12'h15A;
        15'h0711: data = 12'h15E;
        15'h0712: data = 12'h162;
        15'h0713: data = 12'h162;
        15'h0714: data = 12'h167;
        15'h0715: data = 12'h169;
        15'h0716: data = 12'h167;
        15'h0717: data = 12'h169;
        15'h0718: data = 12'h16D;
        15'h0719: data = 12'h16B;
        15'h071A: data = 12'h164;
        15'h071B: data = 12'h160;
        15'h071C: data = 12'h165;
        15'h071D: data = 12'h164;
        15'h071E: data = 12'h163;
        15'h071F: data = 12'h16E;
        15'h0720: data = 12'h16F;
        15'h0721: data = 12'h17B;
        15'h0722: data = 12'h17F;
        15'h0723: data = 12'h18D;
        15'h0724: data = 12'h193;
        15'h0725: data = 12'h196;
        15'h0726: data = 12'h19C;
        15'h0727: data = 12'h1A2;
        15'h0728: data = 12'h1AD;
        15'h0729: data = 12'h1AD;
        15'h072A: data = 12'h1AB;
        15'h072B: data = 12'h1AB;
        15'h072C: data = 12'h1B1;
        15'h072D: data = 12'h1BA;
        15'h072E: data = 12'h1C0;
        15'h072F: data = 12'h1C6;
        15'h0730: data = 12'h1D0;
        15'h0731: data = 12'h1DB;
        15'h0732: data = 12'h1E6;
        15'h0733: data = 12'h1F4;
        15'h0734: data = 12'h205;
        15'h0735: data = 12'h211;
        15'h0736: data = 12'h21A;
        15'h0737: data = 12'h222;
        15'h0738: data = 12'h22E;
        15'h0739: data = 12'h236;
        15'h073A: data = 12'h240;
        15'h073B: data = 12'h24A;
        15'h073C: data = 12'h256;
        15'h073D: data = 12'h257;
        15'h073E: data = 12'h267;
        15'h073F: data = 12'h26C;
        15'h0740: data = 12'h27A;
        15'h0741: data = 12'h282;
        15'h0742: data = 12'h293;
        15'h0743: data = 12'h2A0;
        15'h0744: data = 12'h2B4;
        15'h0745: data = 12'h2C5;
        15'h0746: data = 12'h2D5;
        15'h0747: data = 12'h2E6;
        15'h0748: data = 12'h2FA;
        15'h0749: data = 12'h30B;
        15'h074A: data = 12'h318;
        15'h074B: data = 12'h32A;
        15'h074C: data = 12'h336;
        15'h074D: data = 12'h344;
        15'h074E: data = 12'h352;
        15'h074F: data = 12'h35E;
        15'h0750: data = 12'h36A;
        15'h0751: data = 12'h376;
        15'h0752: data = 12'h389;
        15'h0753: data = 12'h390;
        15'h0754: data = 12'h3A6;
        15'h0755: data = 12'h3B8;
        15'h0756: data = 12'h3C8;
        15'h0757: data = 12'h3DC;
        15'h0758: data = 12'h3F3;
        15'h0759: data = 12'h404;
        15'h075A: data = 12'h419;
        15'h075B: data = 12'h433;
        15'h075C: data = 12'h446;
        15'h075D: data = 12'h45F;
        15'h075E: data = 12'h46E;
        15'h075F: data = 12'h482;
        15'h0760: data = 12'h490;
        15'h0761: data = 12'h4A7;
        15'h0762: data = 12'h4B8;
        15'h0763: data = 12'h4CB;
        15'h0764: data = 12'h4D8;
        15'h0765: data = 12'h4ED;
        15'h0766: data = 12'h501;
        15'h0767: data = 12'h50D;
        15'h0768: data = 12'h523;
        15'h0769: data = 12'h53A;
        15'h076A: data = 12'h54F;
        15'h076B: data = 12'h560;
        15'h076C: data = 12'h573;
        15'h076D: data = 12'h58A;
        15'h076E: data = 12'h5A3;
        15'h076F: data = 12'h5B8;
        15'h0770: data = 12'h5D4;
        15'h0771: data = 12'h5EE;
        15'h0772: data = 12'h604;
        15'h0773: data = 12'h61F;
        15'h0774: data = 12'h631;
        15'h0775: data = 12'h649;
        15'h0776: data = 12'h660;
        15'h0777: data = 12'h676;
        15'h0778: data = 12'h68A;
        15'h0779: data = 12'h69F;
        15'h077A: data = 12'h6B5;
        15'h077B: data = 12'h6C9;
        15'h077C: data = 12'h6DA;
        15'h077D: data = 12'h6ED;
        15'h077E: data = 12'h704;
        15'h077F: data = 12'h719;
        15'h0780: data = 12'h731;
        15'h0781: data = 12'h745;
        15'h0782: data = 12'h758;
        15'h0783: data = 12'h777;
        15'h0784: data = 12'h78C;
        15'h0785: data = 12'h7A6;
        15'h0786: data = 12'h7C1;
        15'h0787: data = 12'h7D9;
        15'h0788: data = 12'h7F1;
        15'h0789: data = 12'h809;
        15'h078A: data = 12'h089;
        15'h078B: data = 12'h08D;
        15'h078C: data = 12'h0A4;
        15'h078D: data = 12'h0B3;
        15'h078E: data = 12'h0CE;
        15'h078F: data = 12'h0E9;
        15'h0790: data = 12'h0FF;
        15'h0791: data = 12'h10D;
        15'h0792: data = 12'h127;
        15'h0793: data = 12'h13C;
        15'h0794: data = 12'h14C;
        15'h0795: data = 12'h161;
        15'h0796: data = 12'h174;
        15'h0797: data = 12'h18B;
        15'h0798: data = 12'h1A8;
        15'h0799: data = 12'h1BA;
        15'h079A: data = 12'h1CF;
        15'h079B: data = 12'h1EC;
        15'h079C: data = 12'h206;
        15'h079D: data = 12'h215;
        15'h079E: data = 12'h22F;
        15'h079F: data = 12'h24F;
        15'h07A0: data = 12'h265;
        15'h07A1: data = 12'h279;
        15'h07A2: data = 12'h292;
        15'h07A3: data = 12'h2AE;
        15'h07A4: data = 12'h2CA;
        15'h07A5: data = 12'h2DC;
        15'h07A6: data = 12'h2FA;
        15'h07A7: data = 12'h30B;
        15'h07A8: data = 12'h326;
        15'h07A9: data = 12'h33B;
        15'h07AA: data = 12'h352;
        15'h07AB: data = 12'h367;
        15'h07AC: data = 12'h37C;
        15'h07AD: data = 12'h398;
        15'h07AE: data = 12'h3A9;
        15'h07AF: data = 12'h3BF;
        15'h07B0: data = 12'h3D6;
        15'h07B1: data = 12'h3EC;
        15'h07B2: data = 12'h3FC;
        15'h07B3: data = 12'h415;
        15'h07B4: data = 12'h428;
        15'h07B5: data = 12'h43C;
        15'h07B6: data = 12'h44A;
        15'h07B7: data = 12'h45F;
        15'h07B8: data = 12'h474;
        15'h07B9: data = 12'h488;
        15'h07BA: data = 12'h49B;
        15'h07BB: data = 12'h4AD;
        15'h07BC: data = 12'h4BE;
        15'h07BD: data = 12'h4D7;
        15'h07BE: data = 12'h4EB;
        15'h07BF: data = 12'h4FF;
        15'h07C0: data = 12'h50A;
        15'h07C1: data = 12'h521;
        15'h07C2: data = 12'h538;
        15'h07C3: data = 12'h546;
        15'h07C4: data = 12'h55F;
        15'h07C5: data = 12'h56E;
        15'h07C6: data = 12'h584;
        15'h07C7: data = 12'h594;
        15'h07C8: data = 12'h5A8;
        15'h07C9: data = 12'h5BF;
        15'h07CA: data = 12'h5CB;
        15'h07CB: data = 12'h5DD;
        15'h07CC: data = 12'h5F3;
        15'h07CD: data = 12'h606;
        15'h07CE: data = 12'h616;
        15'h07CF: data = 12'h628;
        15'h07D0: data = 12'h638;
        15'h07D1: data = 12'h643;
        15'h07D2: data = 12'h656;
        15'h07D3: data = 12'h66D;
        15'h07D4: data = 12'h67A;
        15'h07D5: data = 12'h686;
        15'h07D6: data = 12'h698;
        15'h07D7: data = 12'h6A8;
        15'h07D8: data = 12'h6B5;
        15'h07D9: data = 12'h6C5;
        15'h07DA: data = 12'h6D5;
        15'h07DB: data = 12'h6DE;
        15'h07DC: data = 12'h6F0;
        15'h07DD: data = 12'h700;
        15'h07DE: data = 12'h704;
        15'h07DF: data = 12'h714;
        15'h07E0: data = 12'h724;
        15'h07E1: data = 12'h732;
        15'h07E2: data = 12'h736;
        15'h07E3: data = 12'h73D;
        15'h07E4: data = 12'h74E;
        15'h07E5: data = 12'h760;
        15'h07E6: data = 12'h766;
        15'h07E7: data = 12'h772;
        15'h07E8: data = 12'h779;
        15'h07E9: data = 12'h787;
        15'h07EA: data = 12'h78E;
        15'h07EB: data = 12'h797;
        15'h07EC: data = 12'h79D;
        15'h07ED: data = 12'h7A5;
        15'h07EE: data = 12'h7AE;
        15'h07EF: data = 12'h7B6;
        15'h07F0: data = 12'h7BD;
        15'h07F1: data = 12'h7C2;
        15'h07F2: data = 12'h7CA;
        15'h07F3: data = 12'h7D2;
        15'h07F4: data = 12'h7DC;
        15'h07F5: data = 12'h7E3;
        15'h07F6: data = 12'h7E6;
        15'h07F7: data = 12'h7ED;
        15'h07F8: data = 12'h7F3;
        15'h07F9: data = 12'h7F6;
        15'h07FA: data = 12'h7FC;
        15'h07FB: data = 12'h805;
        15'h07FC: data = 12'h494;
        15'h07FD: data = 12'h083;
        15'h07FE: data = 12'h090;
        15'h07FF: data = 12'h095;
        15'h0800: data = 12'h097;
        15'h0801: data = 12'h0A0;
        15'h0802: data = 12'h0A1;
        15'h0803: data = 12'h0AE;
        15'h0804: data = 12'h0AD;
        15'h0805: data = 12'h0B1;
        15'h0806: data = 12'h0BF;
        15'h0807: data = 12'h0C0;
        15'h0808: data = 12'h0C2;
        15'h0809: data = 12'h0C5;
        15'h080A: data = 12'h0D2;
        15'h080B: data = 12'h0D3;
        15'h080C: data = 12'h0D5;
        15'h080D: data = 12'h0D4;
        15'h080E: data = 12'h0D8;
        15'h080F: data = 12'h0D3;
        15'h0810: data = 12'h0D1;
        15'h0811: data = 12'h0C8;
        15'h0812: data = 12'h0C7;
        15'h0813: data = 12'h0C2;
        15'h0814: data = 12'h0BE;
        15'h0815: data = 12'h0BD;
        15'h0816: data = 12'h0B2;
        15'h0817: data = 12'h0B4;
        15'h0818: data = 12'h0AF;
        15'h0819: data = 12'h0B3;
        15'h081A: data = 12'h0AF;
        15'h081B: data = 12'h0B2;
        15'h081C: data = 12'h0B5;
        15'h081D: data = 12'h0B5;
        15'h081E: data = 12'h0AD;
        15'h081F: data = 12'h0A8;
        15'h0820: data = 12'h0A0;
        15'h0821: data = 12'h091;
        15'h0822: data = 12'h087;
        15'h0823: data = 12'h07B;
        15'h0824: data = 12'h075;
        15'h0825: data = 12'h079;
        15'h0826: data = 12'h079;
        15'h0827: data = 12'h078;
        15'h0828: data = 12'h06D;
        15'h0829: data = 12'h065;
        15'h082A: data = 12'h05C;
        15'h082B: data = 12'h050;
        15'h082C: data = 12'h042;
        15'h082D: data = 12'h02E;
        15'h082E: data = 12'h7B3;
        15'h082F: data = 12'h7AC;
        15'h0830: data = 12'h7AE;
        15'h0831: data = 12'h7A5;
        15'h0832: data = 12'h798;
        15'h0833: data = 12'h78F;
        15'h0834: data = 12'h777;
        15'h0835: data = 12'h768;
        15'h0836: data = 12'h752;
        15'h0837: data = 12'h74A;
        15'h0838: data = 12'h73C;
        15'h0839: data = 12'h739;
        15'h083A: data = 12'h730;
        15'h083B: data = 12'h726;
        15'h083C: data = 12'h71C;
        15'h083D: data = 12'h70B;
        15'h083E: data = 12'h6F5;
        15'h083F: data = 12'h6E0;
        15'h0840: data = 12'h6D1;
        15'h0841: data = 12'h6BF;
        15'h0842: data = 12'h6B1;
        15'h0843: data = 12'h6AA;
        15'h0844: data = 12'h69E;
        15'h0845: data = 12'h68F;
        15'h0846: data = 12'h688;
        15'h0847: data = 12'h678;
        15'h0848: data = 12'h668;
        15'h0849: data = 12'h658;
        15'h084A: data = 12'h642;
        15'h084B: data = 12'h62F;
        15'h084C: data = 12'h61D;
        15'h084D: data = 12'h605;
        15'h084E: data = 12'h5F8;
        15'h084F: data = 12'h5E7;
        15'h0850: data = 12'h5D8;
        15'h0851: data = 12'h5C6;
        15'h0852: data = 12'h5BC;
        15'h0853: data = 12'h5B3;
        15'h0854: data = 12'h59E;
        15'h0855: data = 12'h590;
        15'h0856: data = 12'h575;
        15'h0857: data = 12'h567;
        15'h0858: data = 12'h554;
        15'h0859: data = 12'h53F;
        15'h085A: data = 12'h528;
        15'h085B: data = 12'h512;
        15'h085C: data = 12'h4FE;
        15'h085D: data = 12'h4E5;
        15'h085E: data = 12'h4CC;
        15'h085F: data = 12'h4BC;
        15'h0860: data = 12'h4A7;
        15'h0861: data = 12'h495;
        15'h0862: data = 12'h483;
        15'h0863: data = 12'h46C;
        15'h0864: data = 12'h458;
        15'h0865: data = 12'h44A;
        15'h0866: data = 12'h435;
        15'h0867: data = 12'h420;
        15'h0868: data = 12'h40A;
        15'h0869: data = 12'h3F7;
        15'h086A: data = 12'h3E9;
        15'h086B: data = 12'h3D6;
        15'h086C: data = 12'h3BC;
        15'h086D: data = 12'h3A3;
        15'h086E: data = 12'h390;
        15'h086F: data = 12'h37A;
        15'h0870: data = 12'h360;
        15'h0871: data = 12'h34A;
        15'h0872: data = 12'h339;
        15'h0873: data = 12'h324;
        15'h0874: data = 12'h308;
        15'h0875: data = 12'h2F1;
        15'h0876: data = 12'h2DB;
        15'h0877: data = 12'h2C3;
        15'h0878: data = 12'h2AC;
        15'h0879: data = 12'h292;
        15'h087A: data = 12'h27C;
        15'h087B: data = 12'h265;
        15'h087C: data = 12'h24A;
        15'h087D: data = 12'h237;
        15'h087E: data = 12'h21B;
        15'h087F: data = 12'h208;
        15'h0880: data = 12'h1F3;
        15'h0881: data = 12'h1D5;
        15'h0882: data = 12'h1BB;
        15'h0883: data = 12'h1A2;
        15'h0884: data = 12'h18F;
        15'h0885: data = 12'h179;
        15'h0886: data = 12'h15B;
        15'h0887: data = 12'h146;
        15'h0888: data = 12'h12F;
        15'h0889: data = 12'h119;
        15'h088A: data = 12'h0FF;
        15'h088B: data = 12'h0E9;
        15'h088C: data = 12'h0D4;
        15'h088D: data = 12'h0BC;
        15'h088E: data = 12'h09D;
        15'h088F: data = 12'h08B;
        15'h0890: data = 12'h077;
        15'h0891: data = 12'h05A;
        15'h0892: data = 12'h041;
        15'h0893: data = 12'h7DB;
        15'h0894: data = 12'h7C7;
        15'h0895: data = 12'h7AD;
        15'h0896: data = 12'h797;
        15'h0897: data = 12'h780;
        15'h0898: data = 12'h76C;
        15'h0899: data = 12'h752;
        15'h089A: data = 12'h740;
        15'h089B: data = 12'h725;
        15'h089C: data = 12'h70C;
        15'h089D: data = 12'h6FA;
        15'h089E: data = 12'h6E1;
        15'h089F: data = 12'h6CB;
        15'h08A0: data = 12'h6B8;
        15'h08A1: data = 12'h69F;
        15'h08A2: data = 12'h686;
        15'h08A3: data = 12'h677;
        15'h08A4: data = 12'h659;
        15'h08A5: data = 12'h64A;
        15'h08A6: data = 12'h62B;
        15'h08A7: data = 12'h619;
        15'h08A8: data = 12'h605;
        15'h08A9: data = 12'h5EE;
        15'h08AA: data = 12'h5DA;
        15'h08AB: data = 12'h5C4;
        15'h08AC: data = 12'h5B1;
        15'h08AD: data = 12'h597;
        15'h08AE: data = 12'h580;
        15'h08AF: data = 12'h56D;
        15'h08B0: data = 12'h55E;
        15'h08B1: data = 12'h551;
        15'h08B2: data = 12'h539;
        15'h08B3: data = 12'h522;
        15'h08B4: data = 12'h512;
        15'h08B5: data = 12'h4FF;
        15'h08B6: data = 12'h4EB;
        15'h08B7: data = 12'h4DE;
        15'h08B8: data = 12'h4C6;
        15'h08B9: data = 12'h4B9;
        15'h08BA: data = 12'h4A1;
        15'h08BB: data = 12'h493;
        15'h08BC: data = 12'h47B;
        15'h08BD: data = 12'h468;
        15'h08BE: data = 12'h457;
        15'h08BF: data = 12'h445;
        15'h08C0: data = 12'h42D;
        15'h08C1: data = 12'h41D;
        15'h08C2: data = 12'h405;
        15'h08C3: data = 12'h3F7;
        15'h08C4: data = 12'h3DE;
        15'h08C5: data = 12'h3CC;
        15'h08C6: data = 12'h3B5;
        15'h08C7: data = 12'h3A3;
        15'h08C8: data = 12'h38F;
        15'h08C9: data = 12'h37F;
        15'h08CA: data = 12'h36C;
        15'h08CB: data = 12'h35C;
        15'h08CC: data = 12'h34F;
        15'h08CD: data = 12'h340;
        15'h08CE: data = 12'h331;
        15'h08CF: data = 12'h32B;
        15'h08D0: data = 12'h31A;
        15'h08D1: data = 12'h30D;
        15'h08D2: data = 12'h301;
        15'h08D3: data = 12'h2F2;
        15'h08D4: data = 12'h2E4;
        15'h08D5: data = 12'h2DA;
        15'h08D6: data = 12'h2C6;
        15'h08D7: data = 12'h2BA;
        15'h08D8: data = 12'h2A7;
        15'h08D9: data = 12'h299;
        15'h08DA: data = 12'h289;
        15'h08DB: data = 12'h273;
        15'h08DC: data = 12'h26C;
        15'h08DD: data = 12'h25C;
        15'h08DE: data = 12'h255;
        15'h08DF: data = 12'h244;
        15'h08E0: data = 12'h23F;
        15'h08E1: data = 12'h234;
        15'h08E2: data = 12'h230;
        15'h08E3: data = 12'h226;
        15'h08E4: data = 12'h222;
        15'h08E5: data = 12'h21A;
        15'h08E6: data = 12'h210;
        15'h08E7: data = 12'h202;
        15'h08E8: data = 12'h1F8;
        15'h08E9: data = 12'h1EE;
        15'h08EA: data = 12'h1E0;
        15'h08EB: data = 12'h1D6;
        15'h08EC: data = 12'h1CA;
        15'h08ED: data = 12'h1BE;
        15'h08EE: data = 12'h1B9;
        15'h08EF: data = 12'h1B1;
        15'h08F0: data = 12'h1AA;
        15'h08F1: data = 12'h1A9;
        15'h08F2: data = 12'h1A2;
        15'h08F3: data = 12'h1A4;
        15'h08F4: data = 12'h1A3;
        15'h08F5: data = 12'h19F;
        15'h08F6: data = 12'h197;
        15'h08F7: data = 12'h195;
        15'h08F8: data = 12'h18D;
        15'h08F9: data = 12'h181;
        15'h08FA: data = 12'h17E;
        15'h08FB: data = 12'h16F;
        15'h08FC: data = 12'h16B;
        15'h08FD: data = 12'h163;
        15'h08FE: data = 12'h164;
        15'h08FF: data = 12'h167;
        15'h0900: data = 12'h161;
        15'h0901: data = 12'h163;
        15'h0902: data = 12'h16A;
        15'h0903: data = 12'h16A;
        15'h0904: data = 12'h165;
        15'h0905: data = 12'h168;
        15'h0906: data = 12'h167;
        15'h0907: data = 12'h166;
        15'h0908: data = 12'h162;
        15'h0909: data = 12'h161;
        15'h090A: data = 12'h15E;
        15'h090B: data = 12'h15C;
        15'h090C: data = 12'h15F;
        15'h090D: data = 12'h15F;
        15'h090E: data = 12'h15D;
        15'h090F: data = 12'h15C;
        15'h0910: data = 12'h16B;
        15'h0911: data = 12'h16C;
        15'h0912: data = 12'h16F;
        15'h0913: data = 12'h17B;
        15'h0914: data = 12'h17D;
        15'h0915: data = 12'h188;
        15'h0916: data = 12'h18B;
        15'h0917: data = 12'h18D;
        15'h0918: data = 12'h193;
        15'h0919: data = 12'h18F;
        15'h091A: data = 12'h193;
        15'h091B: data = 12'h19A;
        15'h091C: data = 12'h19E;
        15'h091D: data = 12'h1A0;
        15'h091E: data = 12'h19F;
        15'h091F: data = 12'h1AC;
        15'h0920: data = 12'h1B1;
        15'h0921: data = 12'h1BC;
        15'h0922: data = 12'h1C5;
        15'h0923: data = 12'h1D3;
        15'h0924: data = 12'h1DD;
        15'h0925: data = 12'h1E7;
        15'h0926: data = 12'h1F1;
        15'h0927: data = 12'h1FA;
        15'h0928: data = 12'h208;
        15'h0929: data = 12'h20D;
        15'h092A: data = 12'h216;
        15'h092B: data = 12'h21A;
        15'h092C: data = 12'h222;
        15'h092D: data = 12'h228;
        15'h092E: data = 12'h232;
        15'h092F: data = 12'h23B;
        15'h0930: data = 12'h247;
        15'h0931: data = 12'h252;
        15'h0932: data = 12'h262;
        15'h0933: data = 12'h26D;
        15'h0934: data = 12'h284;
        15'h0935: data = 12'h28B;
        15'h0936: data = 12'h29E;
        15'h0937: data = 12'h2B2;
        15'h0938: data = 12'h2C0;
        15'h0939: data = 12'h2D1;
        15'h093A: data = 12'h2DA;
        15'h093B: data = 12'h2E8;
        15'h093C: data = 12'h2F8;
        15'h093D: data = 12'h303;
        15'h093E: data = 12'h310;
        15'h093F: data = 12'h31C;
        15'h0940: data = 12'h32C;
        15'h0941: data = 12'h332;
        15'h0942: data = 12'h341;
        15'h0943: data = 12'h353;
        15'h0944: data = 12'h362;
        15'h0945: data = 12'h36F;
        15'h0946: data = 12'h38A;
        15'h0947: data = 12'h394;
        15'h0948: data = 12'h3AC;
        15'h0949: data = 12'h3C5;
        15'h094A: data = 12'h3D5;
        15'h094B: data = 12'h3EC;
        15'h094C: data = 12'h400;
        15'h094D: data = 12'h411;
        15'h094E: data = 12'h426;
        15'h094F: data = 12'h433;
        15'h0950: data = 12'h445;
        15'h0951: data = 12'h45A;
        15'h0952: data = 12'h463;
        15'h0953: data = 12'h47A;
        15'h0954: data = 12'h489;
        15'h0955: data = 12'h49D;
        15'h0956: data = 12'h4A9;
        15'h0957: data = 12'h4BF;
        15'h0958: data = 12'h4CA;
        15'h0959: data = 12'h4E4;
        15'h095A: data = 12'h4FA;
        15'h095B: data = 12'h50C;
        15'h095C: data = 12'h525;
        15'h095D: data = 12'h53C;
        15'h095E: data = 12'h556;
        15'h095F: data = 12'h56D;
        15'h0960: data = 12'h581;
        15'h0961: data = 12'h59C;
        15'h0962: data = 12'h5AF;
        15'h0963: data = 12'h5C5;
        15'h0964: data = 12'h5DC;
        15'h0965: data = 12'h5F1;
        15'h0966: data = 12'h605;
        15'h0967: data = 12'h620;
        15'h0968: data = 12'h62C;
        15'h0969: data = 12'h63F;
        15'h096A: data = 12'h655;
        15'h096B: data = 12'h664;
        15'h096C: data = 12'h682;
        15'h096D: data = 12'h68E;
        15'h096E: data = 12'h6A6;
        15'h096F: data = 12'h6BD;
        15'h0970: data = 12'h6D3;
        15'h0971: data = 12'h6E9;
        15'h0972: data = 12'h703;
        15'h0973: data = 12'h71B;
        15'h0974: data = 12'h733;
        15'h0975: data = 12'h74C;
        15'h0976: data = 12'h765;
        15'h0977: data = 12'h780;
        15'h0978: data = 12'h79B;
        15'h0979: data = 12'h7AF;
        15'h097A: data = 12'h7CA;
        15'h097B: data = 12'h7E0;
        15'h097C: data = 12'h7F4;
        15'h097D: data = 12'h80D;
        15'h097E: data = 12'h06C;
        15'h097F: data = 12'h08A;
        15'h0980: data = 12'h0A0;
        15'h0981: data = 12'h0AD;
        15'h0982: data = 12'h0C5;
        15'h0983: data = 12'h0DC;
        15'h0984: data = 12'h0ED;
        15'h0985: data = 12'h0FF;
        15'h0986: data = 12'h114;
        15'h0987: data = 12'h12D;
        15'h0988: data = 12'h144;
        15'h0989: data = 12'h15D;
        15'h098A: data = 12'h171;
        15'h098B: data = 12'h18E;
        15'h098C: data = 12'h1AA;
        15'h098D: data = 12'h1BC;
        15'h098E: data = 12'h1DD;
        15'h098F: data = 12'h1F5;
        15'h0990: data = 12'h213;
        15'h0991: data = 12'h223;
        15'h0992: data = 12'h240;
        15'h0993: data = 12'h25C;
        15'h0994: data = 12'h271;
        15'h0995: data = 12'h286;
        15'h0996: data = 12'h29B;
        15'h0997: data = 12'h2B6;
        15'h0998: data = 12'h2CE;
        15'h0999: data = 12'h2DC;
        15'h099A: data = 12'h2F7;
        15'h099B: data = 12'h309;
        15'h099C: data = 12'h326;
        15'h099D: data = 12'h336;
        15'h099E: data = 12'h34A;
        15'h099F: data = 12'h360;
        15'h09A0: data = 12'h373;
        15'h09A1: data = 12'h389;
        15'h09A2: data = 12'h39E;
        15'h09A3: data = 12'h3B6;
        15'h09A4: data = 12'h3C8;
        15'h09A5: data = 12'h3DC;
        15'h09A6: data = 12'h3F0;
        15'h09A7: data = 12'h409;
        15'h09A8: data = 12'h41F;
        15'h09A9: data = 12'h436;
        15'h09AA: data = 12'h446;
        15'h09AB: data = 12'h459;
        15'h09AC: data = 12'h472;
        15'h09AD: data = 12'h485;
        15'h09AE: data = 12'h49C;
        15'h09AF: data = 12'h4B2;
        15'h09B0: data = 12'h4C2;
        15'h09B1: data = 12'h4DC;
        15'h09B2: data = 12'h4F1;
        15'h09B3: data = 12'h508;
        15'h09B4: data = 12'h515;
        15'h09B5: data = 12'h52E;
        15'h09B6: data = 12'h547;
        15'h09B7: data = 12'h551;
        15'h09B8: data = 12'h569;
        15'h09B9: data = 12'h57B;
        15'h09BA: data = 12'h594;
        15'h09BB: data = 12'h5A5;
        15'h09BC: data = 12'h5B5;
        15'h09BD: data = 12'h5CA;
        15'h09BE: data = 12'h5D7;
        15'h09BF: data = 12'h5E6;
        15'h09C0: data = 12'h5FA;
        15'h09C1: data = 12'h60E;
        15'h09C2: data = 12'h61D;
        15'h09C3: data = 12'h62C;
        15'h09C4: data = 12'h63D;
        15'h09C5: data = 12'h647;
        15'h09C6: data = 12'h65A;
        15'h09C7: data = 12'h66D;
        15'h09C8: data = 12'h67D;
        15'h09C9: data = 12'h685;
        15'h09CA: data = 12'h69A;
        15'h09CB: data = 12'h6A3;
        15'h09CC: data = 12'h6B3;
        15'h09CD: data = 12'h6C6;
        15'h09CE: data = 12'h6D2;
        15'h09CF: data = 12'h6D7;
        15'h09D0: data = 12'h6E7;
        15'h09D1: data = 12'h6F7;
        15'h09D2: data = 12'h6FF;
        15'h09D3: data = 12'h70C;
        15'h09D4: data = 12'h719;
        15'h09D5: data = 12'h723;
        15'h09D6: data = 12'h72C;
        15'h09D7: data = 12'h733;
        15'h09D8: data = 12'h742;
        15'h09D9: data = 12'h750;
        15'h09DA: data = 12'h754;
        15'h09DB: data = 12'h769;
        15'h09DC: data = 12'h770;
        15'h09DD: data = 12'h77B;
        15'h09DE: data = 12'h785;
        15'h09DF: data = 12'h78C;
        15'h09E0: data = 12'h794;
        15'h09E1: data = 12'h79F;
        15'h09E2: data = 12'h7A6;
        15'h09E3: data = 12'h7AE;
        15'h09E4: data = 12'h7B8;
        15'h09E5: data = 12'h7C1;
        15'h09E6: data = 12'h7C8;
        15'h09E7: data = 12'h7CE;
        15'h09E8: data = 12'h7DC;
        15'h09E9: data = 12'h7E2;
        15'h09EA: data = 12'h7EA;
        15'h09EB: data = 12'h7F2;
        15'h09EC: data = 12'h7FC;
        15'h09ED: data = 12'h7FE;
        15'h09EE: data = 12'h806;
        15'h09EF: data = 12'h272;
        15'h09F0: data = 12'h08F;
        15'h09F1: data = 12'h090;
        15'h09F2: data = 12'h09D;
        15'h09F3: data = 12'h0A3;
        15'h09F4: data = 12'h0A6;
        15'h09F5: data = 12'h0AE;
        15'h09F6: data = 12'h0B5;
        15'h09F7: data = 12'h0BD;
        15'h09F8: data = 12'h0BE;
        15'h09F9: data = 12'h0BD;
        15'h09FA: data = 12'h0CA;
        15'h09FB: data = 12'h0C9;
        15'h09FC: data = 12'h0CA;
        15'h09FD: data = 12'h0C8;
        15'h09FE: data = 12'h0D3;
        15'h09FF: data = 12'h0D1;
        15'h0A00: data = 12'h0CF;
        15'h0A01: data = 12'h0CB;
        15'h0A02: data = 12'h0C7;
        15'h0A03: data = 12'h0C5;
        15'h0A04: data = 12'h0C5;
        15'h0A05: data = 12'h0BA;
        15'h0A06: data = 12'h0BD;
        15'h0A07: data = 12'h0BF;
        15'h0A08: data = 12'h0C0;
        15'h0A09: data = 12'h0C3;
        15'h0A0A: data = 12'h0C2;
        15'h0A0B: data = 12'h0C7;
        15'h0A0C: data = 12'h0BD;
        15'h0A0D: data = 12'h0BF;
        15'h0A0E: data = 12'h0B9;
        15'h0A0F: data = 12'h0B6;
        15'h0A10: data = 12'h0B3;
        15'h0A11: data = 12'h0AD;
        15'h0A12: data = 12'h09F;
        15'h0A13: data = 12'h097;
        15'h0A14: data = 12'h090;
        15'h0A15: data = 12'h08C;
        15'h0A16: data = 12'h089;
        15'h0A17: data = 12'h08B;
        15'h0A18: data = 12'h088;
        15'h0A19: data = 12'h088;
        15'h0A1A: data = 12'h07E;
        15'h0A1B: data = 12'h075;
        15'h0A1C: data = 12'h068;
        15'h0A1D: data = 12'h05B;
        15'h0A1E: data = 12'h04F;
        15'h0A1F: data = 12'h04A;
        15'h0A20: data = 12'h043;
        15'h0A21: data = 12'h000;
        15'h0A22: data = 12'h7C9;
        15'h0A23: data = 12'h7BD;
        15'h0A24: data = 12'h7B2;
        15'h0A25: data = 12'h7A1;
        15'h0A26: data = 12'h78B;
        15'h0A27: data = 12'h77E;
        15'h0A28: data = 12'h76E;
        15'h0A29: data = 12'h764;
        15'h0A2A: data = 12'h75D;
        15'h0A2B: data = 12'h754;
        15'h0A2C: data = 12'h748;
        15'h0A2D: data = 12'h741;
        15'h0A2E: data = 12'h72F;
        15'h0A2F: data = 12'h724;
        15'h0A30: data = 12'h70A;
        15'h0A31: data = 12'h6FB;
        15'h0A32: data = 12'h6E9;
        15'h0A33: data = 12'h6DD;
        15'h0A34: data = 12'h6D9;
        15'h0A35: data = 12'h6D1;
        15'h0A36: data = 12'h6C4;
        15'h0A37: data = 12'h6B9;
        15'h0A38: data = 12'h6A8;
        15'h0A39: data = 12'h695;
        15'h0A3A: data = 12'h67F;
        15'h0A3B: data = 12'h66B;
        15'h0A3C: data = 12'h656;
        15'h0A3D: data = 12'h646;
        15'h0A3E: data = 12'h636;
        15'h0A3F: data = 12'h626;
        15'h0A40: data = 12'h623;
        15'h0A41: data = 12'h615;
        15'h0A42: data = 12'h607;
        15'h0A43: data = 12'h5F6;
        15'h0A44: data = 12'h5E3;
        15'h0A45: data = 12'h5D1;
        15'h0A46: data = 12'h5C1;
        15'h0A47: data = 12'h5B1;
        15'h0A48: data = 12'h595;
        15'h0A49: data = 12'h584;
        15'h0A4A: data = 12'h566;
        15'h0A4B: data = 12'h556;
        15'h0A4C: data = 12'h545;
        15'h0A4D: data = 12'h533;
        15'h0A4E: data = 12'h51C;
        15'h0A4F: data = 12'h50B;
        15'h0A50: data = 12'h4FE;
        15'h0A51: data = 12'h4EB;
        15'h0A52: data = 12'h4D5;
        15'h0A53: data = 12'h4C7;
        15'h0A54: data = 12'h4B8;
        15'h0A55: data = 12'h4A6;
        15'h0A56: data = 12'h493;
        15'h0A57: data = 12'h47F;
        15'h0A58: data = 12'h468;
        15'h0A59: data = 12'h454;
        15'h0A5A: data = 12'h43F;
        15'h0A5B: data = 12'h427;
        15'h0A5C: data = 12'h40D;
        15'h0A5D: data = 12'h3F9;
        15'h0A5E: data = 12'h3E4;
        15'h0A5F: data = 12'h3CF;
        15'h0A60: data = 12'h3B5;
        15'h0A61: data = 12'h3A0;
        15'h0A62: data = 12'h388;
        15'h0A63: data = 12'h36B;
        15'h0A64: data = 12'h353;
        15'h0A65: data = 12'h33D;
        15'h0A66: data = 12'h32C;
        15'h0A67: data = 12'h315;
        15'h0A68: data = 12'h2F7;
        15'h0A69: data = 12'h2E3;
        15'h0A6A: data = 12'h2CD;
        15'h0A6B: data = 12'h2B8;
        15'h0A6C: data = 12'h29C;
        15'h0A6D: data = 12'h281;
        15'h0A6E: data = 12'h26E;
        15'h0A6F: data = 12'h256;
        15'h0A70: data = 12'h23C;
        15'h0A71: data = 12'h228;
        15'h0A72: data = 12'h20F;
        15'h0A73: data = 12'h1FB;
        15'h0A74: data = 12'h1E8;
        15'h0A75: data = 12'h1CB;
        15'h0A76: data = 12'h1B3;
        15'h0A77: data = 12'h199;
        15'h0A78: data = 12'h185;
        15'h0A79: data = 12'h169;
        15'h0A7A: data = 12'h153;
        15'h0A7B: data = 12'h13C;
        15'h0A7C: data = 12'h127;
        15'h0A7D: data = 12'h10F;
        15'h0A7E: data = 12'h0FB;
        15'h0A7F: data = 12'h0E3;
        15'h0A80: data = 12'h0CE;
        15'h0A81: data = 12'h0B4;
        15'h0A82: data = 12'h098;
        15'h0A83: data = 12'h083;
        15'h0A84: data = 12'h070;
        15'h0A85: data = 12'h055;
        15'h0A86: data = 12'h03E;
        15'h0A87: data = 12'h7CD;
        15'h0A88: data = 12'h7BE;
        15'h0A89: data = 12'h7A8;
        15'h0A8A: data = 12'h795;
        15'h0A8B: data = 12'h77B;
        15'h0A8C: data = 12'h764;
        15'h0A8D: data = 12'h74F;
        15'h0A8E: data = 12'h73B;
        15'h0A8F: data = 12'h725;
        15'h0A90: data = 12'h70F;
        15'h0A91: data = 12'h6F7;
        15'h0A92: data = 12'h6E1;
        15'h0A93: data = 12'h6CC;
        15'h0A94: data = 12'h6B9;
        15'h0A95: data = 12'h6A0;
        15'h0A96: data = 12'h689;
        15'h0A97: data = 12'h67A;
        15'h0A98: data = 12'h65F;
        15'h0A99: data = 12'h64E;
        15'h0A9A: data = 12'h635;
        15'h0A9B: data = 12'h625;
        15'h0A9C: data = 12'h60E;
        15'h0A9D: data = 12'h5FA;
        15'h0A9E: data = 12'h5E4;
        15'h0A9F: data = 12'h5D0;
        15'h0AA0: data = 12'h5BF;
        15'h0AA1: data = 12'h5A8;
        15'h0AA2: data = 12'h593;
        15'h0AA3: data = 12'h57F;
        15'h0AA4: data = 12'h56C;
        15'h0AA5: data = 12'h55A;
        15'h0AA6: data = 12'h545;
        15'h0AA7: data = 12'h52D;
        15'h0AA8: data = 12'h51C;
        15'h0AA9: data = 12'h508;
        15'h0AAA: data = 12'h4F0;
        15'h0AAB: data = 12'h4DD;
        15'h0AAC: data = 12'h4C6;
        15'h0AAD: data = 12'h4B4;
        15'h0AAE: data = 12'h49D;
        15'h0AAF: data = 12'h48B;
        15'h0AB0: data = 12'h477;
        15'h0AB1: data = 12'h45D;
        15'h0AB2: data = 12'h44A;
        15'h0AB3: data = 12'h438;
        15'h0AB4: data = 12'h41E;
        15'h0AB5: data = 12'h40D;
        15'h0AB6: data = 12'h3F6;
        15'h0AB7: data = 12'h3E4;
        15'h0AB8: data = 12'h3D6;
        15'h0AB9: data = 12'h3C3;
        15'h0ABA: data = 12'h3B0;
        15'h0ABB: data = 12'h3A1;
        15'h0ABC: data = 12'h391;
        15'h0ABD: data = 12'h389;
        15'h0ABE: data = 12'h378;
        15'h0ABF: data = 12'h36B;
        15'h0AC0: data = 12'h35D;
        15'h0AC1: data = 12'h34D;
        15'h0AC2: data = 12'h340;
        15'h0AC3: data = 12'h330;
        15'h0AC4: data = 12'h31F;
        15'h0AC5: data = 12'h30E;
        15'h0AC6: data = 12'h2FE;
        15'h0AC7: data = 12'h2ED;
        15'h0AC8: data = 12'h2DA;
        15'h0AC9: data = 12'h2D0;
        15'h0ACA: data = 12'h2BB;
        15'h0ACB: data = 12'h2AB;
        15'h0ACC: data = 12'h29C;
        15'h0ACD: data = 12'h291;
        15'h0ACE: data = 12'h284;
        15'h0ACF: data = 12'h272;
        15'h0AD0: data = 12'h270;
        15'h0AD1: data = 12'h263;
        15'h0AD2: data = 12'h25E;
        15'h0AD3: data = 12'h252;
        15'h0AD4: data = 12'h24E;
        15'h0AD5: data = 12'h23C;
        15'h0AD6: data = 12'h236;
        15'h0AD7: data = 12'h229;
        15'h0AD8: data = 12'h21E;
        15'h0AD9: data = 12'h216;
        15'h0ADA: data = 12'h208;
        15'h0ADB: data = 12'h1F7;
        15'h0ADC: data = 12'h1E7;
        15'h0ADD: data = 12'h1E0;
        15'h0ADE: data = 12'h1DA;
        15'h0ADF: data = 12'h1D1;
        15'h0AE0: data = 12'h1CA;
        15'h0AE1: data = 12'h1C1;
        15'h0AE2: data = 12'h1C0;
        15'h0AE3: data = 12'h1BD;
        15'h0AE4: data = 12'h1BA;
        15'h0AE5: data = 12'h1B5;
        15'h0AE6: data = 12'h1A8;
        15'h0AE7: data = 12'h1A9;
        15'h0AE8: data = 12'h1A3;
        15'h0AE9: data = 12'h197;
        15'h0AEA: data = 12'h18C;
        15'h0AEB: data = 12'h188;
        15'h0AEC: data = 12'h17D;
        15'h0AED: data = 12'h173;
        15'h0AEE: data = 12'h173;
        15'h0AEF: data = 12'h16C;
        15'h0AF0: data = 12'h171;
        15'h0AF1: data = 12'h16C;
        15'h0AF2: data = 12'h16E;
        15'h0AF3: data = 12'h175;
        15'h0AF4: data = 12'h170;
        15'h0AF5: data = 12'h170;
        15'h0AF6: data = 12'h170;
        15'h0AF7: data = 12'h16F;
        15'h0AF8: data = 12'h164;
        15'h0AF9: data = 12'h15E;
        15'h0AFA: data = 12'h15F;
        15'h0AFB: data = 12'h156;
        15'h0AFC: data = 12'h155;
        15'h0AFD: data = 12'h157;
        15'h0AFE: data = 12'h156;
        15'h0AFF: data = 12'h15D;
        15'h0B00: data = 12'h161;
        15'h0B01: data = 12'h164;
        15'h0B02: data = 12'h166;
        15'h0B03: data = 12'h16C;
        15'h0B04: data = 12'h178;
        15'h0B05: data = 12'h178;
        15'h0B06: data = 12'h177;
        15'h0B07: data = 12'h17D;
        15'h0B08: data = 12'h17C;
        15'h0B09: data = 12'h180;
        15'h0B0A: data = 12'h182;
        15'h0B0B: data = 12'h17E;
        15'h0B0C: data = 12'h183;
        15'h0B0D: data = 12'h183;
        15'h0B0E: data = 12'h18B;
        15'h0B0F: data = 12'h195;
        15'h0B10: data = 12'h19B;
        15'h0B11: data = 12'h1A6;
        15'h0B12: data = 12'h1AA;
        15'h0B13: data = 12'h1B8;
        15'h0B14: data = 12'h1C2;
        15'h0B15: data = 12'h1CD;
        15'h0B16: data = 12'h1D4;
        15'h0B17: data = 12'h1DB;
        15'h0B18: data = 12'h1E1;
        15'h0B19: data = 12'h1E8;
        15'h0B1A: data = 12'h1ED;
        15'h0B1B: data = 12'h1F4;
        15'h0B1C: data = 12'h1FB;
        15'h0B1D: data = 12'h201;
        15'h0B1E: data = 12'h209;
        15'h0B1F: data = 12'h20F;
        15'h0B20: data = 12'h21F;
        15'h0B21: data = 12'h221;
        15'h0B22: data = 12'h234;
        15'h0B23: data = 12'h243;
        15'h0B24: data = 12'h255;
        15'h0B25: data = 12'h261;
        15'h0B26: data = 12'h272;
        15'h0B27: data = 12'h27C;
        15'h0B28: data = 12'h28C;
        15'h0B29: data = 12'h293;
        15'h0B2A: data = 12'h2A5;
        15'h0B2B: data = 12'h2B3;
        15'h0B2C: data = 12'h2BE;
        15'h0B2D: data = 12'h2C8;
        15'h0B2E: data = 12'h2CE;
        15'h0B2F: data = 12'h2DA;
        15'h0B30: data = 12'h2EA;
        15'h0B31: data = 12'h2F7;
        15'h0B32: data = 12'h308;
        15'h0B33: data = 12'h317;
        15'h0B34: data = 12'h328;
        15'h0B35: data = 12'h335;
        15'h0B36: data = 12'h34A;
        15'h0B37: data = 12'h35E;
        15'h0B38: data = 12'h371;
        15'h0B39: data = 12'h384;
        15'h0B3A: data = 12'h39A;
        15'h0B3B: data = 12'h3A3;
        15'h0B3C: data = 12'h3B7;
        15'h0B3D: data = 12'h3C9;
        15'h0B3E: data = 12'h3D6;
        15'h0B3F: data = 12'h3EC;
        15'h0B40: data = 12'h3FB;
        15'h0B41: data = 12'h40C;
        15'h0B42: data = 12'h41A;
        15'h0B43: data = 12'h428;
        15'h0B44: data = 12'h436;
        15'h0B45: data = 12'h44A;
        15'h0B46: data = 12'h459;
        15'h0B47: data = 12'h471;
        15'h0B48: data = 12'h480;
        15'h0B49: data = 12'h498;
        15'h0B4A: data = 12'h4A9;
        15'h0B4B: data = 12'h4C4;
        15'h0B4C: data = 12'h4D8;
        15'h0B4D: data = 12'h4F1;
        15'h0B4E: data = 12'h50C;
        15'h0B4F: data = 12'h51C;
        15'h0B50: data = 12'h532;
        15'h0B51: data = 12'h54B;
        15'h0B52: data = 12'h55F;
        15'h0B53: data = 12'h572;
        15'h0B54: data = 12'h583;
        15'h0B55: data = 12'h594;
        15'h0B56: data = 12'h5A9;
        15'h0B57: data = 12'h5BB;
        15'h0B58: data = 12'h5D4;
        15'h0B59: data = 12'h5E7;
        15'h0B5A: data = 12'h5F8;
        15'h0B5B: data = 12'h60F;
        15'h0B5C: data = 12'h622;
        15'h0B5D: data = 12'h636;
        15'h0B5E: data = 12'h64A;
        15'h0B5F: data = 12'h665;
        15'h0B60: data = 12'h682;
        15'h0B61: data = 12'h695;
        15'h0B62: data = 12'h6AE;
        15'h0B63: data = 12'h6C8;
        15'h0B64: data = 12'h6E1;
        15'h0B65: data = 12'h6F7;
        15'h0B66: data = 12'h714;
        15'h0B67: data = 12'h72A;
        15'h0B68: data = 12'h741;
        15'h0B69: data = 12'h757;
        15'h0B6A: data = 12'h76C;
        15'h0B6B: data = 12'h780;
        15'h0B6C: data = 12'h79B;
        15'h0B6D: data = 12'h7AD;
        15'h0B6E: data = 12'h7C4;
        15'h0B6F: data = 12'h7D7;
        15'h0B70: data = 12'h7EB;
        15'h0B71: data = 12'h7FD;
        15'h0B72: data = 12'h066;
        15'h0B73: data = 12'h07E;
        15'h0B74: data = 12'h092;
        15'h0B75: data = 12'h0A0;
        15'h0B76: data = 12'h0BD;
        15'h0B77: data = 12'h0D6;
        15'h0B78: data = 12'h0F1;
        15'h0B79: data = 12'h102;
        15'h0B7A: data = 12'h121;
        15'h0B7B: data = 12'h136;
        15'h0B7C: data = 12'h153;
        15'h0B7D: data = 12'h16A;
        15'h0B7E: data = 12'h183;
        15'h0B7F: data = 12'h19D;
        15'h0B80: data = 12'h1B8;
        15'h0B81: data = 12'h1C8;
        15'h0B82: data = 12'h1E4;
        15'h0B83: data = 12'h1FC;
        15'h0B84: data = 12'h212;
        15'h0B85: data = 12'h223;
        15'h0B86: data = 12'h240;
        15'h0B87: data = 12'h256;
        15'h0B88: data = 12'h26D;
        15'h0B89: data = 12'h27E;
        15'h0B8A: data = 12'h28E;
        15'h0B8B: data = 12'h2A8;
        15'h0B8C: data = 12'h2C2;
        15'h0B8D: data = 12'h2D2;
        15'h0B8E: data = 12'h2E9;
        15'h0B8F: data = 12'h2FF;
        15'h0B90: data = 12'h316;
        15'h0B91: data = 12'h329;
        15'h0B92: data = 12'h33F;
        15'h0B93: data = 12'h357;
        15'h0B94: data = 12'h36C;
        15'h0B95: data = 12'h386;
        15'h0B96: data = 12'h39B;
        15'h0B97: data = 12'h3B3;
        15'h0B98: data = 12'h3CD;
        15'h0B99: data = 12'h3E2;
        15'h0B9A: data = 12'h3F7;
        15'h0B9B: data = 12'h40E;
        15'h0B9C: data = 12'h426;
        15'h0B9D: data = 12'h43E;
        15'h0B9E: data = 12'h452;
        15'h0B9F: data = 12'h467;
        15'h0BA0: data = 12'h480;
        15'h0BA1: data = 12'h497;
        15'h0BA2: data = 12'h4A9;
        15'h0BA3: data = 12'h4C2;
        15'h0BA4: data = 12'h4D1;
        15'h0BA5: data = 12'h4E9;
        15'h0BA6: data = 12'h4FE;
        15'h0BA7: data = 12'h512;
        15'h0BA8: data = 12'h51D;
        15'h0BA9: data = 12'h535;
        15'h0BAA: data = 12'h54D;
        15'h0BAB: data = 12'h556;
        15'h0BAC: data = 12'h56B;
        15'h0BAD: data = 12'h57D;
        15'h0BAE: data = 12'h591;
        15'h0BAF: data = 12'h5A2;
        15'h0BB0: data = 12'h5B3;
        15'h0BB1: data = 12'h5C9;
        15'h0BB2: data = 12'h5D4;
        15'h0BB3: data = 12'h5E1;
        15'h0BB4: data = 12'h5F5;
        15'h0BB5: data = 12'h608;
        15'h0BB6: data = 12'h614;
        15'h0BB7: data = 12'h623;
        15'h0BB8: data = 12'h631;
        15'h0BB9: data = 12'h63B;
        15'h0BBA: data = 12'h64C;
        15'h0BBB: data = 12'h65F;
        15'h0BBC: data = 12'h670;
        15'h0BBD: data = 12'h679;
        15'h0BBE: data = 12'h68E;
        15'h0BBF: data = 12'h697;
        15'h0BC0: data = 12'h6A5;
        15'h0BC1: data = 12'h6B5;
        15'h0BC2: data = 12'h6C3;
        15'h0BC3: data = 12'h6CE;
        15'h0BC4: data = 12'h6DF;
        15'h0BC5: data = 12'h6EC;
        15'h0BC6: data = 12'h6F4;
        15'h0BC7: data = 12'h702;
        15'h0BC8: data = 12'h713;
        15'h0BC9: data = 12'h722;
        15'h0BCA: data = 12'h729;
        15'h0BCB: data = 12'h733;
        15'h0BCC: data = 12'h740;
        15'h0BCD: data = 12'h74F;
        15'h0BCE: data = 12'h758;
        15'h0BCF: data = 12'h76B;
        15'h0BD0: data = 12'h770;
        15'h0BD1: data = 12'h77F;
        15'h0BD2: data = 12'h78A;
        15'h0BD3: data = 12'h790;
        15'h0BD4: data = 12'h79B;
        15'h0BD5: data = 12'h7A7;
        15'h0BD6: data = 12'h7B4;
        15'h0BD7: data = 12'h7BF;
        15'h0BD8: data = 12'h7C7;
        15'h0BD9: data = 12'h7CE;
        15'h0BDA: data = 12'h7D5;
        15'h0BDB: data = 12'h7DE;
        15'h0BDC: data = 12'h7E8;
        15'h0BDD: data = 12'h7EE;
        15'h0BDE: data = 12'h7F7;
        15'h0BDF: data = 12'h800;
        15'h0BE0: data = 12'h807;
        15'h0BE1: data = 12'h808;
        15'h0BE2: data = 12'h811;
        15'h0BE3: data = 12'h819;
        15'h0BE4: data = 12'h099;
        15'h0BE5: data = 12'h09B;
        15'h0BE6: data = 12'h0A7;
        15'h0BE7: data = 12'h0A8;
        15'h0BE8: data = 12'h0AB;
        15'h0BE9: data = 12'h0B3;
        15'h0BEA: data = 12'h0B2;
        15'h0BEB: data = 12'h0BD;
        15'h0BEC: data = 12'h0BF;
        15'h0BED: data = 12'h0BC;
        15'h0BEE: data = 12'h0C5;
        15'h0BEF: data = 12'h0C3;
        15'h0BF0: data = 12'h0C0;
        15'h0BF1: data = 12'h0BF;
        15'h0BF2: data = 12'h0C7;
        15'h0BF3: data = 12'h0C6;
        15'h0BF4: data = 12'h0C5;
        15'h0BF5: data = 12'h0C2;
        15'h0BF6: data = 12'h0C1;
        15'h0BF7: data = 12'h0C3;
        15'h0BF8: data = 12'h0C7;
        15'h0BF9: data = 12'h0C0;
        15'h0BFA: data = 12'h0C7;
        15'h0BFB: data = 12'h0CA;
        15'h0BFC: data = 12'h0CB;
        15'h0BFD: data = 12'h0D1;
        15'h0BFE: data = 12'h0C9;
        15'h0BFF: data = 12'h0C9;
        15'h0C00: data = 12'h0BB;
        15'h0C01: data = 12'h0BB;
        15'h0C02: data = 12'h0B0;
        15'h0C03: data = 12'h0AA;
        15'h0C04: data = 12'h0A3;
        15'h0C05: data = 12'h0A2;
        15'h0C06: data = 12'h09C;
        15'h0C07: data = 12'h099;
        15'h0C08: data = 12'h09F;
        15'h0C09: data = 12'h09B;
        15'h0C0A: data = 12'h096;
        15'h0C0B: data = 12'h08E;
        15'h0C0C: data = 12'h086;
        15'h0C0D: data = 12'h084;
        15'h0C0E: data = 12'h076;
        15'h0C0F: data = 12'h067;
        15'h0C10: data = 12'h05E;
        15'h0C11: data = 12'h057;
        15'h0C12: data = 12'h053;
        15'h0C13: data = 12'h056;
        15'h0C14: data = 12'h04E;
        15'h0C15: data = 12'h08D;
        15'h0C16: data = 12'h7C1;
        15'h0C17: data = 12'h7B4;
        15'h0C18: data = 12'h7A2;
        15'h0C19: data = 12'h794;
        15'h0C1A: data = 12'h785;
        15'h0C1B: data = 12'h780;
        15'h0C1C: data = 12'h776;
        15'h0C1D: data = 12'h771;
        15'h0C1E: data = 12'h762;
        15'h0C1F: data = 12'h757;
        15'h0C20: data = 12'h746;
        15'h0C21: data = 12'h739;
        15'h0C22: data = 12'h725;
        15'h0C23: data = 12'h715;
        15'h0C24: data = 12'h708;
        15'h0C25: data = 12'h6FC;
        15'h0C26: data = 12'h6F1;
        15'h0C27: data = 12'h6EA;
        15'h0C28: data = 12'h6E3;
        15'h0C29: data = 12'h6D6;
        15'h0C2A: data = 12'h6C3;
        15'h0C2B: data = 12'h6B2;
        15'h0C2C: data = 12'h69E;
        15'h0C2D: data = 12'h688;
        15'h0C2E: data = 12'h674;
        15'h0C2F: data = 12'h664;
        15'h0C30: data = 12'h658;
        15'h0C31: data = 12'h64C;
        15'h0C32: data = 12'h641;
        15'h0C33: data = 12'h636;
        15'h0C34: data = 12'h62E;
        15'h0C35: data = 12'h618;
        15'h0C36: data = 12'h607;
        15'h0C37: data = 12'h5F6;
        15'h0C38: data = 12'h5DD;
        15'h0C39: data = 12'h5C8;
        15'h0C3A: data = 12'h5B6;
        15'h0C3B: data = 12'h5A4;
        15'h0C3C: data = 12'h58A;
        15'h0C3D: data = 12'h57B;
        15'h0C3E: data = 12'h561;
        15'h0C3F: data = 12'h555;
        15'h0C40: data = 12'h54A;
        15'h0C41: data = 12'h538;
        15'h0C42: data = 12'h527;
        15'h0C43: data = 12'h518;
        15'h0C44: data = 12'h508;
        15'h0C45: data = 12'h4F7;
        15'h0C46: data = 12'h4DF;
        15'h0C47: data = 12'h4CB;
        15'h0C48: data = 12'h4B9;
        15'h0C49: data = 12'h4A2;
        15'h0C4A: data = 12'h48D;
        15'h0C4B: data = 12'h47B;
        15'h0C4C: data = 12'h461;
        15'h0C4D: data = 12'h451;
        15'h0C4E: data = 12'h437;
        15'h0C4F: data = 12'h41B;
        15'h0C50: data = 12'h406;
        15'h0C51: data = 12'h3EA;
        15'h0C52: data = 12'h3D8;
        15'h0C53: data = 12'h3C5;
        15'h0C54: data = 12'h3AB;
        15'h0C55: data = 12'h390;
        15'h0C56: data = 12'h37C;
        15'h0C57: data = 12'h365;
        15'h0C58: data = 12'h34D;
        15'h0C59: data = 12'h337;
        15'h0C5A: data = 12'h323;
        15'h0C5B: data = 12'h311;
        15'h0C5C: data = 12'h2F6;
        15'h0C5D: data = 12'h2E2;
        15'h0C5E: data = 12'h2CB;
        15'h0C5F: data = 12'h2B8;
        15'h0C60: data = 12'h29C;
        15'h0C61: data = 12'h284;
        15'h0C62: data = 12'h274;
        15'h0C63: data = 12'h25D;
        15'h0C64: data = 12'h241;
        15'h0C65: data = 12'h22F;
        15'h0C66: data = 12'h211;
        15'h0C67: data = 12'h1FE;
        15'h0C68: data = 12'h1ED;
        15'h0C69: data = 12'h1D0;
        15'h0C6A: data = 12'h1B8;
        15'h0C6B: data = 12'h19F;
        15'h0C6C: data = 12'h18F;
        15'h0C6D: data = 12'h176;
        15'h0C6E: data = 12'h15D;
        15'h0C6F: data = 12'h145;
        15'h0C70: data = 12'h12F;
        15'h0C71: data = 12'h11A;
        15'h0C72: data = 12'h101;
        15'h0C73: data = 12'h0EC;
        15'h0C74: data = 12'h0D4;
        15'h0C75: data = 12'h0BC;
        15'h0C76: data = 12'h0A2;
        15'h0C77: data = 12'h08E;
        15'h0C78: data = 12'h07C;
        15'h0C79: data = 12'h063;
        15'h0C7A: data = 12'h047;
        15'h0C7B: data = 12'h7E3;
        15'h0C7C: data = 12'h7CA;
        15'h0C7D: data = 12'h7B6;
        15'h0C7E: data = 12'h79F;
        15'h0C7F: data = 12'h787;
        15'h0C80: data = 12'h771;
        15'h0C81: data = 12'h75E;
        15'h0C82: data = 12'h748;
        15'h0C83: data = 12'h732;
        15'h0C84: data = 12'h71D;
        15'h0C85: data = 12'h704;
        15'h0C86: data = 12'h6F0;
        15'h0C87: data = 12'h6D9;
        15'h0C88: data = 12'h6C2;
        15'h0C89: data = 12'h6AB;
        15'h0C8A: data = 12'h696;
        15'h0C8B: data = 12'h686;
        15'h0C8C: data = 12'h66C;
        15'h0C8D: data = 12'h659;
        15'h0C8E: data = 12'h640;
        15'h0C8F: data = 12'h632;
        15'h0C90: data = 12'h616;
        15'h0C91: data = 12'h601;
        15'h0C92: data = 12'h5EB;
        15'h0C93: data = 12'h5D8;
        15'h0C94: data = 12'h5C5;
        15'h0C95: data = 12'h5AA;
        15'h0C96: data = 12'h595;
        15'h0C97: data = 12'h57D;
        15'h0C98: data = 12'h56D;
        15'h0C99: data = 12'h55C;
        15'h0C9A: data = 12'h53F;
        15'h0C9B: data = 12'h52A;
        15'h0C9C: data = 12'h518;
        15'h0C9D: data = 12'h4FD;
        15'h0C9E: data = 12'h4E7;
        15'h0C9F: data = 12'h4D5;
        15'h0CA0: data = 12'h4BE;
        15'h0CA1: data = 12'h4AA;
        15'h0CA2: data = 12'h48F;
        15'h0CA3: data = 12'h47D;
        15'h0CA4: data = 12'h46B;
        15'h0CA5: data = 12'h453;
        15'h0CA6: data = 12'h443;
        15'h0CA7: data = 12'h433;
        15'h0CA8: data = 12'h41D;
        15'h0CA9: data = 12'h40F;
        15'h0CAA: data = 12'h3F7;
        15'h0CAB: data = 12'h3EA;
        15'h0CAC: data = 12'h3DE;
        15'h0CAD: data = 12'h3CD;
        15'h0CAE: data = 12'h3BC;
        15'h0CAF: data = 12'h3B1;
        15'h0CB0: data = 12'h39D;
        15'h0CB1: data = 12'h394;
        15'h0CB2: data = 12'h383;
        15'h0CB3: data = 12'h36F;
        15'h0CB4: data = 12'h35F;
        15'h0CB5: data = 12'h34E;
        15'h0CB6: data = 12'h33D;
        15'h0CB7: data = 12'h32E;
        15'h0CB8: data = 12'h31B;
        15'h0CB9: data = 12'h305;
        15'h0CBA: data = 12'h2F3;
        15'h0CBB: data = 12'h2E0;
        15'h0CBC: data = 12'h2D1;
        15'h0CBD: data = 12'h2C6;
        15'h0CBE: data = 12'h2B9;
        15'h0CBF: data = 12'h2AD;
        15'h0CC0: data = 12'h29D;
        15'h0CC1: data = 12'h299;
        15'h0CC2: data = 12'h290;
        15'h0CC3: data = 12'h284;
        15'h0CC4: data = 12'h27E;
        15'h0CC5: data = 12'h269;
        15'h0CC6: data = 12'h264;
        15'h0CC7: data = 12'h253;
        15'h0CC8: data = 12'h24D;
        15'h0CC9: data = 12'h23A;
        15'h0CCA: data = 12'h233;
        15'h0CCB: data = 12'h21F;
        15'h0CCC: data = 12'h211;
        15'h0CCD: data = 12'h206;
        15'h0CCE: data = 12'h1FE;
        15'h0CCF: data = 12'h1F2;
        15'h0CD0: data = 12'h1E8;
        15'h0CD1: data = 12'h1DF;
        15'h0CD2: data = 12'h1DF;
        15'h0CD3: data = 12'h1DC;
        15'h0CD4: data = 12'h1D7;
        15'h0CD5: data = 12'h1CE;
        15'h0CD6: data = 12'h1C5;
        15'h0CD7: data = 12'h1C4;
        15'h0CD8: data = 12'h1BB;
        15'h0CD9: data = 12'h1B3;
        15'h0CDA: data = 12'h1A8;
        15'h0CDB: data = 12'h1A0;
        15'h0CDC: data = 12'h197;
        15'h0CDD: data = 12'h189;
        15'h0CDE: data = 12'h181;
        15'h0CDF: data = 12'h183;
        15'h0CE0: data = 12'h17B;
        15'h0CE1: data = 12'h176;
        15'h0CE2: data = 12'h179;
        15'h0CE3: data = 12'h179;
        15'h0CE4: data = 12'h17C;
        15'h0CE5: data = 12'h17A;
        15'h0CE6: data = 12'h179;
        15'h0CE7: data = 12'h178;
        15'h0CE8: data = 12'h16F;
        15'h0CE9: data = 12'h16F;
        15'h0CEA: data = 12'h168;
        15'h0CEB: data = 12'h165;
        15'h0CEC: data = 12'h15A;
        15'h0CED: data = 12'h155;
        15'h0CEE: data = 12'h151;
        15'h0CEF: data = 12'h153;
        15'h0CF0: data = 12'h156;
        15'h0CF1: data = 12'h157;
        15'h0CF2: data = 12'h15B;
        15'h0CF3: data = 12'h167;
        15'h0CF4: data = 12'h16E;
        15'h0CF5: data = 12'h170;
        15'h0CF6: data = 12'h170;
        15'h0CF7: data = 12'h16E;
        15'h0CF8: data = 12'h176;
        15'h0CF9: data = 12'h172;
        15'h0CFA: data = 12'h173;
        15'h0CFB: data = 12'h174;
        15'h0CFC: data = 12'h16F;
        15'h0CFD: data = 12'h176;
        15'h0CFE: data = 12'h179;
        15'h0CFF: data = 12'h17C;
        15'h0D00: data = 12'h184;
        15'h0D01: data = 12'h187;
        15'h0D02: data = 12'h194;
        15'h0D03: data = 12'h19D;
        15'h0D04: data = 12'h1A8;
        15'h0D05: data = 12'h1AF;
        15'h0D06: data = 12'h1B3;
        15'h0D07: data = 12'h1BB;
        15'h0D08: data = 12'h1C1;
        15'h0D09: data = 12'h1CB;
        15'h0D0A: data = 12'h1D1;
        15'h0D0B: data = 12'h1D5;
        15'h0D0C: data = 12'h1DB;
        15'h0D0D: data = 12'h1DE;
        15'h0D0E: data = 12'h1DE;
        15'h0D0F: data = 12'h1E9;
        15'h0D10: data = 12'h1F6;
        15'h0D11: data = 12'h1FD;
        15'h0D12: data = 12'h20A;
        15'h0D13: data = 12'h210;
        15'h0D14: data = 12'h227;
        15'h0D15: data = 12'h232;
        15'h0D16: data = 12'h243;
        15'h0D17: data = 12'h24D;
        15'h0D18: data = 12'h25C;
        15'h0D19: data = 12'h267;
        15'h0D1A: data = 12'h275;
        15'h0D1B: data = 12'h27F;
        15'h0D1C: data = 12'h289;
        15'h0D1D: data = 12'h28D;
        15'h0D1E: data = 12'h29A;
        15'h0D1F: data = 12'h2A7;
        15'h0D20: data = 12'h2AF;
        15'h0D21: data = 12'h2B8;
        15'h0D22: data = 12'h2C6;
        15'h0D23: data = 12'h2D6;
        15'h0D24: data = 12'h2E8;
        15'h0D25: data = 12'h2F7;
        15'h0D26: data = 12'h30E;
        15'h0D27: data = 12'h31C;
        15'h0D28: data = 12'h32F;
        15'h0D29: data = 12'h340;
        15'h0D2A: data = 12'h354;
        15'h0D2B: data = 12'h364;
        15'h0D2C: data = 12'h378;
        15'h0D2D: data = 12'h384;
        15'h0D2E: data = 12'h399;
        15'h0D2F: data = 12'h3A0;
        15'h0D30: data = 12'h3B5;
        15'h0D31: data = 12'h3C3;
        15'h0D32: data = 12'h3D0;
        15'h0D33: data = 12'h3E2;
        15'h0D34: data = 12'h3F1;
        15'h0D35: data = 12'h3FB;
        15'h0D36: data = 12'h411;
        15'h0D37: data = 12'h421;
        15'h0D38: data = 12'h432;
        15'h0D39: data = 12'h44A;
        15'h0D3A: data = 12'h45B;
        15'h0D3B: data = 12'h476;
        15'h0D3C: data = 12'h489;
        15'h0D3D: data = 12'h4A2;
        15'h0D3E: data = 12'h4B4;
        15'h0D3F: data = 12'h4CD;
        15'h0D40: data = 12'h4DE;
        15'h0D41: data = 12'h4F5;
        15'h0D42: data = 12'h50D;
        15'h0D43: data = 12'h51B;
        15'h0D44: data = 12'h533;
        15'h0D45: data = 12'h54A;
        15'h0D46: data = 12'h55A;
        15'h0D47: data = 12'h568;
        15'h0D48: data = 12'h57A;
        15'h0D49: data = 12'h58F;
        15'h0D4A: data = 12'h59D;
        15'h0D4B: data = 12'h5B5;
        15'h0D4C: data = 12'h5C9;
        15'h0D4D: data = 12'h5E0;
        15'h0D4E: data = 12'h5F7;
        15'h0D4F: data = 12'h612;
        15'h0D50: data = 12'h620;
        15'h0D51: data = 12'h63B;
        15'h0D52: data = 12'h658;
        15'h0D53: data = 12'h66E;
        15'h0D54: data = 12'h688;
        15'h0D55: data = 12'h6A1;
        15'h0D56: data = 12'h6B7;
        15'h0D57: data = 12'h6CE;
        15'h0D58: data = 12'h6E5;
        15'h0D59: data = 12'h6FA;
        15'h0D5A: data = 12'h712;
        15'h0D5B: data = 12'h72A;
        15'h0D5C: data = 12'h73F;
        15'h0D5D: data = 12'h752;
        15'h0D5E: data = 12'h764;
        15'h0D5F: data = 12'h779;
        15'h0D60: data = 12'h78F;
        15'h0D61: data = 12'h7A2;
        15'h0D62: data = 12'h7B4;
        15'h0D63: data = 12'h7CF;
        15'h0D64: data = 12'h7E5;
        15'h0D65: data = 12'h7FD;
        15'h0D66: data = 12'h067;
        15'h0D67: data = 12'h081;
        15'h0D68: data = 12'h096;
        15'h0D69: data = 12'h0AA;
        15'h0D6A: data = 12'h0C7;
        15'h0D6B: data = 12'h0E2;
        15'h0D6C: data = 12'h0FC;
        15'h0D6D: data = 12'h10D;
        15'h0D6E: data = 12'h12C;
        15'h0D6F: data = 12'h143;
        15'h0D70: data = 12'h15A;
        15'h0D71: data = 12'h16D;
        15'h0D72: data = 12'h188;
        15'h0D73: data = 12'h19E;
        15'h0D74: data = 12'h1B6;
        15'h0D75: data = 12'h1CB;
        15'h0D76: data = 12'h1DD;
        15'h0D77: data = 12'h1F9;
        15'h0D78: data = 12'h210;
        15'h0D79: data = 12'h21D;
        15'h0D7A: data = 12'h235;
        15'h0D7B: data = 12'h24C;
        15'h0D7C: data = 12'h260;
        15'h0D7D: data = 12'h275;
        15'h0D7E: data = 12'h28A;
        15'h0D7F: data = 12'h2A2;
        15'h0D80: data = 12'h2B9;
        15'h0D81: data = 12'h2C8;
        15'h0D82: data = 12'h2E6;
        15'h0D83: data = 12'h2FA;
        15'h0D84: data = 12'h31A;
        15'h0D85: data = 12'h32B;
        15'h0D86: data = 12'h341;
        15'h0D87: data = 12'h359;
        15'h0D88: data = 12'h375;
        15'h0D89: data = 12'h38F;
        15'h0D8A: data = 12'h3A6;
        15'h0D8B: data = 12'h3C1;
        15'h0D8C: data = 12'h3DA;
        15'h0D8D: data = 12'h3ED;
        15'h0D8E: data = 12'h400;
        15'h0D8F: data = 12'h419;
        15'h0D90: data = 12'h430;
        15'h0D91: data = 12'h444;
        15'h0D92: data = 12'h457;
        15'h0D93: data = 12'h46C;
        15'h0D94: data = 12'h485;
        15'h0D95: data = 12'h496;
        15'h0D96: data = 12'h4AF;
        15'h0D97: data = 12'h4BE;
        15'h0D98: data = 12'h4D0;
        15'h0D99: data = 12'h4E5;
        15'h0D9A: data = 12'h4F8;
        15'h0D9B: data = 12'h50D;
        15'h0D9C: data = 12'h51B;
        15'h0D9D: data = 12'h52D;
        15'h0D9E: data = 12'h541;
        15'h0D9F: data = 12'h551;
        15'h0DA0: data = 12'h564;
        15'h0DA1: data = 12'h56D;
        15'h0DA2: data = 12'h584;
        15'h0DA3: data = 12'h594;
        15'h0DA4: data = 12'h5A4;
        15'h0DA5: data = 12'h5BB;
        15'h0DA6: data = 12'h5C8;
        15'h0DA7: data = 12'h5D5;
        15'h0DA8: data = 12'h5EE;
        15'h0DA9: data = 12'h5FA;
        15'h0DAA: data = 12'h609;
        15'h0DAB: data = 12'h61B;
        15'h0DAC: data = 12'h62A;
        15'h0DAD: data = 12'h636;
        15'h0DAE: data = 12'h649;
        15'h0DAF: data = 12'h65D;
        15'h0DB0: data = 12'h66D;
        15'h0DB1: data = 12'h679;
        15'h0DB2: data = 12'h68C;
        15'h0DB3: data = 12'h699;
        15'h0DB4: data = 12'h6A8;
        15'h0DB5: data = 12'h6BA;
        15'h0DB6: data = 12'h6C5;
        15'h0DB7: data = 12'h6D3;
        15'h0DB8: data = 12'h6E5;
        15'h0DB9: data = 12'h6F6;
        15'h0DBA: data = 12'h6FD;
        15'h0DBB: data = 12'h70C;
        15'h0DBC: data = 12'h71D;
        15'h0DBD: data = 12'h72F;
        15'h0DBE: data = 12'h733;
        15'h0DBF: data = 12'h73E;
        15'h0DC0: data = 12'h74D;
        15'h0DC1: data = 12'h760;
        15'h0DC2: data = 12'h767;
        15'h0DC3: data = 12'h777;
        15'h0DC4: data = 12'h77E;
        15'h0DC5: data = 12'h78D;
        15'h0DC6: data = 12'h796;
        15'h0DC7: data = 12'h7A2;
        15'h0DC8: data = 12'h7A7;
        15'h0DC9: data = 12'h7B0;
        15'h0DCA: data = 12'h7B8;
        15'h0DCB: data = 12'h7C4;
        15'h0DCC: data = 12'h7CB;
        15'h0DCD: data = 12'h7D1;
        15'h0DCE: data = 12'h7D6;
        15'h0DCF: data = 12'h7E5;
        15'h0DD0: data = 12'h7E7;
        15'h0DD1: data = 12'h7EF;
        15'h0DD2: data = 12'h7F4;
        15'h0DD3: data = 12'h7FE;
        15'h0DD4: data = 12'h802;
        15'h0DD5: data = 12'h803;
        15'h0DD6: data = 12'h80C;
        15'h0DD7: data = 12'h814;
        15'h0DD8: data = 12'h8A2;
        15'h0DD9: data = 12'h093;
        15'h0DDA: data = 12'h09D;
        15'h0DDB: data = 12'h0A1;
        15'h0DDC: data = 12'h0A0;
        15'h0DDD: data = 12'h0A6;
        15'h0DDE: data = 12'h0A5;
        15'h0DDF: data = 12'h0AD;
        15'h0DE0: data = 12'h0AF;
        15'h0DE1: data = 12'h0AD;
        15'h0DE2: data = 12'h0B8;
        15'h0DE3: data = 12'h0B5;
        15'h0DE4: data = 12'h0B7;
        15'h0DE5: data = 12'h0B8;
        15'h0DE6: data = 12'h0C1;
        15'h0DE7: data = 12'h0C3;
        15'h0DE8: data = 12'h0C7;
        15'h0DE9: data = 12'h0C5;
        15'h0DEA: data = 12'h0C9;
        15'h0DEB: data = 12'h0CB;
        15'h0DEC: data = 12'h0CF;
        15'h0DED: data = 12'h0CC;
        15'h0DEE: data = 12'h0CC;
        15'h0DEF: data = 12'h0CE;
        15'h0DF0: data = 12'h0CE;
        15'h0DF1: data = 12'h0CA;
        15'h0DF2: data = 12'h0C6;
        15'h0DF3: data = 12'h0C0;
        15'h0DF4: data = 12'h0B2;
        15'h0DF5: data = 12'h0B1;
        15'h0DF6: data = 12'h0AA;
        15'h0DF7: data = 12'h0A1;
        15'h0DF8: data = 12'h0A5;
        15'h0DF9: data = 12'h0A7;
        15'h0DFA: data = 12'h0A3;
        15'h0DFB: data = 12'h09E;
        15'h0DFC: data = 12'h0A4;
        15'h0DFD: data = 12'h09D;
        15'h0DFE: data = 12'h094;
        15'h0DFF: data = 12'h08A;
        15'h0E00: data = 12'h07F;
        15'h0E01: data = 12'h079;
        15'h0E02: data = 12'h06C;
        15'h0E03: data = 12'h063;
        15'h0E04: data = 12'h05E;
        15'h0E05: data = 12'h05B;
        15'h0E06: data = 12'h05C;
        15'h0E07: data = 12'h058;
        15'h0E08: data = 12'h04C;
        15'h0E09: data = 12'h03C;
        15'h0E0A: data = 12'h7C0;
        15'h0E0B: data = 12'h7AD;
        15'h0E0C: data = 12'h79E;
        15'h0E0D: data = 12'h790;
        15'h0E0E: data = 12'h78A;
        15'h0E0F: data = 12'h785;
        15'h0E10: data = 12'h77C;
        15'h0E11: data = 12'h775;
        15'h0E12: data = 12'h760;
        15'h0E13: data = 12'h755;
        15'h0E14: data = 12'h73C;
        15'h0E15: data = 12'h732;
        15'h0E16: data = 12'h721;
        15'h0E17: data = 12'h716;
        15'h0E18: data = 12'h70C;
        15'h0E19: data = 12'h707;
        15'h0E1A: data = 12'h6F9;
        15'h0E1B: data = 12'h6ED;
        15'h0E1C: data = 12'h6E4;
        15'h0E1D: data = 12'h6D3;
        15'h0E1E: data = 12'h6BE;
        15'h0E1F: data = 12'h6AD;
        15'h0E20: data = 12'h695;
        15'h0E21: data = 12'h687;
        15'h0E22: data = 12'h675;
        15'h0E23: data = 12'h664;
        15'h0E24: data = 12'h65C;
        15'h0E25: data = 12'h654;
        15'h0E26: data = 12'h647;
        15'h0E27: data = 12'h639;
        15'h0E28: data = 12'h631;
        15'h0E29: data = 12'h617;
        15'h0E2A: data = 12'h606;
        15'h0E2B: data = 12'h5EE;
        15'h0E2C: data = 12'h5D8;
        15'h0E2D: data = 12'h5C1;
        15'h0E2E: data = 12'h5AE;
        15'h0E2F: data = 12'h5A2;
        15'h0E30: data = 12'h58C;
        15'h0E31: data = 12'h57E;
        15'h0E32: data = 12'h568;
        15'h0E33: data = 12'h55C;
        15'h0E34: data = 12'h552;
        15'h0E35: data = 12'h541;
        15'h0E36: data = 12'h530;
        15'h0E37: data = 12'h51C;
        15'h0E38: data = 12'h50B;
        15'h0E39: data = 12'h4F5;
        15'h0E3A: data = 12'h4DE;
        15'h0E3B: data = 12'h4CA;
        15'h0E3C: data = 12'h4B7;
        15'h0E3D: data = 12'h4A2;
        15'h0E3E: data = 12'h48C;
        15'h0E3F: data = 12'h475;
        15'h0E40: data = 12'h45D;
        15'h0E41: data = 12'h448;
        15'h0E42: data = 12'h431;
        15'h0E43: data = 12'h415;
        15'h0E44: data = 12'h3FE;
        15'h0E45: data = 12'h3E9;
        15'h0E46: data = 12'h3D3;
        15'h0E47: data = 12'h3C0;
        15'h0E48: data = 12'h3A6;
        15'h0E49: data = 12'h38F;
        15'h0E4A: data = 12'h37E;
        15'h0E4B: data = 12'h365;
        15'h0E4C: data = 12'h350;
        15'h0E4D: data = 12'h33D;
        15'h0E4E: data = 12'h32A;
        15'h0E4F: data = 12'h315;
        15'h0E50: data = 12'h2F9;
        15'h0E51: data = 12'h2E8;
        15'h0E52: data = 12'h2D0;
        15'h0E53: data = 12'h2BB;
        15'h0E54: data = 12'h2A7;
        15'h0E55: data = 12'h28C;
        15'h0E56: data = 12'h279;
        15'h0E57: data = 12'h266;
        15'h0E58: data = 12'h24A;
        15'h0E59: data = 12'h235;
        15'h0E5A: data = 12'h21A;
        15'h0E5B: data = 12'h207;
        15'h0E5C: data = 12'h1F3;
        15'h0E5D: data = 12'h1D7;
        15'h0E5E: data = 12'h1BF;
        15'h0E5F: data = 12'h1A7;
        15'h0E60: data = 12'h194;
        15'h0E61: data = 12'h17F;
        15'h0E62: data = 12'h165;
        15'h0E63: data = 12'h150;
        15'h0E64: data = 12'h13A;
        15'h0E65: data = 12'h11F;
        15'h0E66: data = 12'h10A;
        15'h0E67: data = 12'h0F6;
        15'h0E68: data = 12'h0DB;
        15'h0E69: data = 12'h0C4;
        15'h0E6A: data = 12'h0A7;
        15'h0E6B: data = 12'h092;
        15'h0E6C: data = 12'h082;
        15'h0E6D: data = 12'h067;
        15'h0E6E: data = 12'h04F;
        15'h0E6F: data = 12'h7E5;
        15'h0E70: data = 12'h7D1;
        15'h0E71: data = 12'h7BC;
        15'h0E72: data = 12'h7A4;
        15'h0E73: data = 12'h790;
        15'h0E74: data = 12'h778;
        15'h0E75: data = 12'h760;
        15'h0E76: data = 12'h74E;
        15'h0E77: data = 12'h735;
        15'h0E78: data = 12'h722;
        15'h0E79: data = 12'h70A;
        15'h0E7A: data = 12'h6F1;
        15'h0E7B: data = 12'h6DB;
        15'h0E7C: data = 12'h6C4;
        15'h0E7D: data = 12'h6AF;
        15'h0E7E: data = 12'h699;
        15'h0E7F: data = 12'h687;
        15'h0E80: data = 12'h66D;
        15'h0E81: data = 12'h659;
        15'h0E82: data = 12'h63F;
        15'h0E83: data = 12'h62E;
        15'h0E84: data = 12'h615;
        15'h0E85: data = 12'h600;
        15'h0E86: data = 12'h5E7;
        15'h0E87: data = 12'h5D2;
        15'h0E88: data = 12'h5C1;
        15'h0E89: data = 12'h5A7;
        15'h0E8A: data = 12'h592;
        15'h0E8B: data = 12'h57A;
        15'h0E8C: data = 12'h568;
        15'h0E8D: data = 12'h552;
        15'h0E8E: data = 12'h53B;
        15'h0E8F: data = 12'h524;
        15'h0E90: data = 12'h512;
        15'h0E91: data = 12'h4F9;
        15'h0E92: data = 12'h4E3;
        15'h0E93: data = 12'h4CF;
        15'h0E94: data = 12'h4B5;
        15'h0E95: data = 12'h4A8;
        15'h0E96: data = 12'h491;
        15'h0E97: data = 12'h47E;
        15'h0E98: data = 12'h46A;
        15'h0E99: data = 12'h455;
        15'h0E9A: data = 12'h447;
        15'h0E9B: data = 12'h43B;
        15'h0E9C: data = 12'h423;
        15'h0E9D: data = 12'h416;
        15'h0E9E: data = 12'h401;
        15'h0E9F: data = 12'h3F5;
        15'h0EA0: data = 12'h3E4;
        15'h0EA1: data = 12'h3D4;
        15'h0EA2: data = 12'h3C0;
        15'h0EA3: data = 12'h3B6;
        15'h0EA4: data = 12'h3A0;
        15'h0EA5: data = 12'h397;
        15'h0EA6: data = 12'h37F;
        15'h0EA7: data = 12'h36D;
        15'h0EA8: data = 12'h35C;
        15'h0EA9: data = 12'h34A;
        15'h0EAA: data = 12'h337;
        15'h0EAB: data = 12'h324;
        15'h0EAC: data = 12'h30F;
        15'h0EAD: data = 12'h2FE;
        15'h0EAE: data = 12'h2EB;
        15'h0EAF: data = 12'h2DB;
        15'h0EB0: data = 12'h2D2;
        15'h0EB1: data = 12'h2CA;
        15'h0EB2: data = 12'h2BE;
        15'h0EB3: data = 12'h2B5;
        15'h0EB4: data = 12'h2A8;
        15'h0EB5: data = 12'h2A1;
        15'h0EB6: data = 12'h298;
        15'h0EB7: data = 12'h282;
        15'h0EB8: data = 12'h27E;
        15'h0EB9: data = 12'h26E;
        15'h0EBA: data = 12'h261;
        15'h0EBB: data = 12'h252;
        15'h0EBC: data = 12'h249;
        15'h0EBD: data = 12'h232;
        15'h0EBE: data = 12'h228;
        15'h0EBF: data = 12'h219;
        15'h0EC0: data = 12'h20E;
        15'h0EC1: data = 12'h209;
        15'h0EC2: data = 12'h201;
        15'h0EC3: data = 12'h1F4;
        15'h0EC4: data = 12'h1ED;
        15'h0EC5: data = 12'h1E9;
        15'h0EC6: data = 12'h1E7;
        15'h0EC7: data = 12'h1E2;
        15'h0EC8: data = 12'h1DE;
        15'h0EC9: data = 12'h1CE;
        15'h0ECA: data = 12'h1C7;
        15'h0ECB: data = 12'h1C4;
        15'h0ECC: data = 12'h1B8;
        15'h0ECD: data = 12'h1AD;
        15'h0ECE: data = 12'h1A0;
        15'h0ECF: data = 12'h197;
        15'h0ED0: data = 12'h194;
        15'h0ED1: data = 12'h18B;
        15'h0ED2: data = 12'h185;
        15'h0ED3: data = 12'h184;
        15'h0ED4: data = 12'h182;
        15'h0ED5: data = 12'h17E;
        15'h0ED6: data = 12'h184;
        15'h0ED7: data = 12'h17D;
        15'h0ED8: data = 12'h17F;
        15'h0ED9: data = 12'h178;
        15'h0EDA: data = 12'h178;
        15'h0EDB: data = 12'h177;
        15'h0EDC: data = 12'h16C;
        15'h0EDD: data = 12'h168;
        15'h0EDE: data = 12'h160;
        15'h0EDF: data = 12'h160;
        15'h0EE0: data = 12'h155;
        15'h0EE1: data = 12'h157;
        15'h0EE2: data = 12'h156;
        15'h0EE3: data = 12'h15A;
        15'h0EE4: data = 12'h160;
        15'h0EE5: data = 12'h166;
        15'h0EE6: data = 12'h166;
        15'h0EE7: data = 12'h16D;
        15'h0EE8: data = 12'h16F;
        15'h0EE9: data = 12'h171;
        15'h0EEA: data = 12'h16D;
        15'h0EEB: data = 12'h16E;
        15'h0EEC: data = 12'h172;
        15'h0EED: data = 12'h170;
        15'h0EEE: data = 12'h169;
        15'h0EEF: data = 12'h171;
        15'h0EF0: data = 12'h16F;
        15'h0EF1: data = 12'h175;
        15'h0EF2: data = 12'h178;
        15'h0EF3: data = 12'h17E;
        15'h0EF4: data = 12'h186;
        15'h0EF5: data = 12'h18A;
        15'h0EF6: data = 12'h197;
        15'h0EF7: data = 12'h1A2;
        15'h0EF8: data = 12'h1AC;
        15'h0EF9: data = 12'h1B2;
        15'h0EFA: data = 12'h1B3;
        15'h0EFB: data = 12'h1BC;
        15'h0EFC: data = 12'h1C0;
        15'h0EFD: data = 12'h1C9;
        15'h0EFE: data = 12'h1CA;
        15'h0EFF: data = 12'h1CC;
        15'h0F00: data = 12'h1D2;
        15'h0F01: data = 12'h1D9;
        15'h0F02: data = 12'h1E1;
        15'h0F03: data = 12'h1E8;
        15'h0F04: data = 12'h1FB;
        15'h0F05: data = 12'h203;
        15'h0F06: data = 12'h210;
        15'h0F07: data = 12'h219;
        15'h0F08: data = 12'h22F;
        15'h0F09: data = 12'h235;
        15'h0F0A: data = 12'h246;
        15'h0F0B: data = 12'h24D;
        15'h0F0C: data = 12'h25C;
        15'h0F0D: data = 12'h263;
        15'h0F0E: data = 12'h274;
        15'h0F0F: data = 12'h27C;
        15'h0F10: data = 12'h285;
        15'h0F11: data = 12'h289;
        15'h0F12: data = 12'h294;
        15'h0F13: data = 12'h2A3;
        15'h0F14: data = 12'h2AD;
        15'h0F15: data = 12'h2BD;
        15'h0F16: data = 12'h2CC;
        15'h0F17: data = 12'h2D9;
        15'h0F18: data = 12'h2EB;
        15'h0F19: data = 12'h2FC;
        15'h0F1A: data = 12'h310;
        15'h0F1B: data = 12'h324;
        15'h0F1C: data = 12'h336;
        15'h0F1D: data = 12'h342;
        15'h0F1E: data = 12'h357;
        15'h0F1F: data = 12'h365;
        15'h0F20: data = 12'h374;
        15'h0F21: data = 12'h382;
        15'h0F22: data = 12'h396;
        15'h0F23: data = 12'h39E;
        15'h0F24: data = 12'h3B3;
        15'h0F25: data = 12'h3BF;
        15'h0F26: data = 12'h3CB;
        15'h0F27: data = 12'h3DD;
        15'h0F28: data = 12'h3ED;
        15'h0F29: data = 12'h3FB;
        15'h0F2A: data = 12'h412;
        15'h0F2B: data = 12'h424;
        15'h0F2C: data = 12'h436;
        15'h0F2D: data = 12'h44C;
        15'h0F2E: data = 12'h463;
        15'h0F2F: data = 12'h47A;
        15'h0F30: data = 12'h48F;
        15'h0F31: data = 12'h4A7;
        15'h0F32: data = 12'h4B8;
        15'h0F33: data = 12'h4D3;
        15'h0F34: data = 12'h4E1;
        15'h0F35: data = 12'h4F6;
        15'h0F36: data = 12'h50A;
        15'h0F37: data = 12'h51B;
        15'h0F38: data = 12'h52C;
        15'h0F39: data = 12'h546;
        15'h0F3A: data = 12'h557;
        15'h0F3B: data = 12'h566;
        15'h0F3C: data = 12'h576;
        15'h0F3D: data = 12'h58C;
        15'h0F3E: data = 12'h59D;
        15'h0F3F: data = 12'h5B0;
        15'h0F40: data = 12'h5CC;
        15'h0F41: data = 12'h5E4;
        15'h0F42: data = 12'h5F9;
        15'h0F43: data = 12'h613;
        15'h0F44: data = 12'h624;
        15'h0F45: data = 12'h63D;
        15'h0F46: data = 12'h65A;
        15'h0F47: data = 12'h66E;
        15'h0F48: data = 12'h68D;
        15'h0F49: data = 12'h69F;
        15'h0F4A: data = 12'h6BA;
        15'h0F4B: data = 12'h6CF;
        15'h0F4C: data = 12'h6E3;
        15'h0F4D: data = 12'h6F9;
        15'h0F4E: data = 12'h712;
        15'h0F4F: data = 12'h727;
        15'h0F50: data = 12'h73D;
        15'h0F51: data = 12'h74C;
        15'h0F52: data = 12'h761;
        15'h0F53: data = 12'h775;
        15'h0F54: data = 12'h78A;
        15'h0F55: data = 12'h79F;
        15'h0F56: data = 12'h7B6;
        15'h0F57: data = 12'h7CC;
        15'h0F58: data = 12'h7E6;
        15'h0F59: data = 12'h7FF;
        15'h0F5A: data = 12'h068;
        15'h0F5B: data = 12'h081;
        15'h0F5C: data = 12'h09C;
        15'h0F5D: data = 12'h0AB;
        15'h0F5E: data = 12'h0C8;
        15'h0F5F: data = 12'h0E7;
        15'h0F60: data = 12'h0FD;
        15'h0F61: data = 12'h10D;
        15'h0F62: data = 12'h12A;
        15'h0F63: data = 12'h142;
        15'h0F64: data = 12'h15C;
        15'h0F65: data = 12'h170;
        15'h0F66: data = 12'h185;
        15'h0F67: data = 12'h19F;
        15'h0F68: data = 12'h1B7;
        15'h0F69: data = 12'h1C7;
        15'h0F6A: data = 12'h1DC;
        15'h0F6B: data = 12'h1F7;
        15'h0F6C: data = 12'h20B;
        15'h0F6D: data = 12'h21A;
        15'h0F6E: data = 12'h235;
        15'h0F6F: data = 12'h24A;
        15'h0F70: data = 12'h25E;
        15'h0F71: data = 12'h273;
        15'h0F72: data = 12'h28A;
        15'h0F73: data = 12'h2A4;
        15'h0F74: data = 12'h2BC;
        15'h0F75: data = 12'h2CC;
        15'h0F76: data = 12'h2E7;
        15'h0F77: data = 12'h2FC;
        15'h0F78: data = 12'h31A;
        15'h0F79: data = 12'h32D;
        15'h0F7A: data = 12'h345;
        15'h0F7B: data = 12'h360;
        15'h0F7C: data = 12'h377;
        15'h0F7D: data = 12'h391;
        15'h0F7E: data = 12'h3A8;
        15'h0F7F: data = 12'h3C1;
        15'h0F80: data = 12'h3DB;
        15'h0F81: data = 12'h3ED;
        15'h0F82: data = 12'h3FD;
        15'h0F83: data = 12'h415;
        15'h0F84: data = 12'h430;
        15'h0F85: data = 12'h446;
        15'h0F86: data = 12'h452;
        15'h0F87: data = 12'h46E;
        15'h0F88: data = 12'h483;
        15'h0F89: data = 12'h498;
        15'h0F8A: data = 12'h4A8;
        15'h0F8B: data = 12'h4BB;
        15'h0F8C: data = 12'h4CD;
        15'h0F8D: data = 12'h4E1;
        15'h0F8E: data = 12'h4F7;
        15'h0F8F: data = 12'h50B;
        15'h0F90: data = 12'h515;
        15'h0F91: data = 12'h52C;
        15'h0F92: data = 12'h541;
        15'h0F93: data = 12'h54A;
        15'h0F94: data = 12'h55F;
        15'h0F95: data = 12'h56C;
        15'h0F96: data = 12'h584;
        15'h0F97: data = 12'h597;
        15'h0F98: data = 12'h5A2;
        15'h0F99: data = 12'h5B9;
        15'h0F9A: data = 12'h5C6;
        15'h0F9B: data = 12'h5D3;
        15'h0F9C: data = 12'h5E8;
        15'h0F9D: data = 12'h5FB;
        15'h0F9E: data = 12'h60B;
        15'h0F9F: data = 12'h619;
        15'h0FA0: data = 12'h62B;
        15'h0FA1: data = 12'h638;
        15'h0FA2: data = 12'h647;
        15'h0FA3: data = 12'h65E;
        15'h0FA4: data = 12'h670;
        15'h0FA5: data = 12'h678;
        15'h0FA6: data = 12'h68D;
        15'h0FA7: data = 12'h69A;
        15'h0FA8: data = 12'h6A8;
        15'h0FA9: data = 12'h6BD;
        15'h0FAA: data = 12'h6C7;
        15'h0FAB: data = 12'h6D9;
        15'h0FAC: data = 12'h6E5;
        15'h0FAD: data = 12'h6F9;
        15'h0FAE: data = 12'h700;
        15'h0FAF: data = 12'h70D;
        15'h0FB0: data = 12'h71F;
        15'h0FB1: data = 12'h730;
        15'h0FB2: data = 12'h735;
        15'h0FB3: data = 12'h73E;
        15'h0FB4: data = 12'h74D;
        15'h0FB5: data = 12'h75D;
        15'h0FB6: data = 12'h767;
        15'h0FB7: data = 12'h775;
        15'h0FB8: data = 12'h77F;
        15'h0FB9: data = 12'h78F;
        15'h0FBA: data = 12'h794;
        15'h0FBB: data = 12'h79D;
        15'h0FBC: data = 12'h7A6;
        15'h0FBD: data = 12'h7B0;
        15'h0FBE: data = 12'h7B7;
        15'h0FBF: data = 12'h7C1;
        15'h0FC0: data = 12'h7CB;
        15'h0FC1: data = 12'h7D1;
        15'h0FC2: data = 12'h7D7;
        15'h0FC3: data = 12'h7E0;
        15'h0FC4: data = 12'h7E5;
        15'h0FC5: data = 12'h7ED;
        15'h0FC6: data = 12'h7F2;
        15'h0FC7: data = 12'h7FC;
        15'h0FC8: data = 12'h802;
        15'h0FC9: data = 12'h803;
        15'h0FCA: data = 12'h80D;
        15'h0FCB: data = 12'h813;
        15'h0FCC: data = 12'h85C;
        15'h0FCD: data = 12'h08F;
        15'h0FCE: data = 12'h09B;
        15'h0FCF: data = 12'h09D;
        15'h0FD0: data = 12'h0A2;
        15'h0FD1: data = 12'h0A5;
        15'h0FD2: data = 12'h0A5;
        15'h0FD3: data = 12'h0AC;
        15'h0FD4: data = 12'h0AE;
        15'h0FD5: data = 12'h0AA;
        15'h0FD6: data = 12'h0B7;
        15'h0FD7: data = 12'h0B7;
        15'h0FD8: data = 12'h0B9;
        15'h0FD9: data = 12'h0B9;
        15'h0FDA: data = 12'h0C0;
        15'h0FDB: data = 12'h0C1;
        15'h0FDC: data = 12'h0C5;
        15'h0FDD: data = 12'h0C7;
        15'h0FDE: data = 12'h0CB;
        15'h0FDF: data = 12'h0CC;
        15'h0FE0: data = 12'h0CF;
        15'h0FE1: data = 12'h0CB;
        15'h0FE2: data = 12'h0CD;
        15'h0FE3: data = 12'h0CD;
        15'h0FE4: data = 12'h0CF;
        15'h0FE5: data = 12'h0CE;
        15'h0FE6: data = 12'h0C3;
        15'h0FE7: data = 12'h0BE;
        15'h0FE8: data = 12'h0B4;
        15'h0FE9: data = 12'h0B2;
        15'h0FEA: data = 12'h0A9;
        15'h0FEB: data = 12'h0A6;
        15'h0FEC: data = 12'h0A6;
        15'h0FED: data = 12'h0AA;
        15'h0FEE: data = 12'h0A5;
        15'h0FEF: data = 12'h0A6;
        15'h0FF0: data = 12'h0A6;
        15'h0FF1: data = 12'h09D;
        15'h0FF2: data = 12'h096;
        15'h0FF3: data = 12'h08A;
        15'h0FF4: data = 12'h080;
        15'h0FF5: data = 12'h079;
        15'h0FF6: data = 12'h06F;
        15'h0FF7: data = 12'h066;
        15'h0FF8: data = 12'h05F;
        15'h0FF9: data = 12'h061;
        15'h0FFA: data = 12'h05F;
        15'h0FFB: data = 12'h058;
        15'h0FFC: data = 12'h04E;
        15'h0FFD: data = 12'h7CA;
        15'h0FFE: data = 12'h7BB;
        15'h0FFF: data = 12'h7AC;
        15'h1000: data = 12'h79D;
        15'h1001: data = 12'h790;
        15'h1002: data = 12'h78A;
        15'h1003: data = 12'h789;
        15'h1004: data = 12'h77B;
        15'h1005: data = 12'h773;
        15'h1006: data = 12'h75F;
        15'h1007: data = 12'h759;
        15'h1008: data = 12'h73C;
        15'h1009: data = 12'h730;
        15'h100A: data = 12'h722;
        15'h100B: data = 12'h714;
        15'h100C: data = 12'h709;
        15'h100D: data = 12'h706;
        15'h100E: data = 12'h6FA;
        15'h100F: data = 12'h6ED;
        15'h1010: data = 12'h6E5;
        15'h1011: data = 12'h6D6;
        15'h1012: data = 12'h6C1;
        15'h1013: data = 12'h6AE;
        15'h1014: data = 12'h696;
        15'h1015: data = 12'h687;
        15'h1016: data = 12'h672;
        15'h1017: data = 12'h668;
        15'h1018: data = 12'h65B;
        15'h1019: data = 12'h652;
        15'h101A: data = 12'h646;
        15'h101B: data = 12'h637;
        15'h101C: data = 12'h62C;
        15'h101D: data = 12'h615;
        15'h101E: data = 12'h604;
        15'h101F: data = 12'h5F4;
        15'h1020: data = 12'h5D6;
        15'h1021: data = 12'h5C3;
        15'h1022: data = 12'h5B3;
        15'h1023: data = 12'h5A1;
        15'h1024: data = 12'h58A;
        15'h1025: data = 12'h57A;
        15'h1026: data = 12'h565;
        15'h1027: data = 12'h559;
        15'h1028: data = 12'h54B;
        15'h1029: data = 12'h53C;
        15'h102A: data = 12'h527;
        15'h102B: data = 12'h51D;
        15'h102C: data = 12'h50A;
        15'h102D: data = 12'h4F7;
        15'h102E: data = 12'h4DB;
        15'h102F: data = 12'h4CD;
        15'h1030: data = 12'h4B9;
        15'h1031: data = 12'h4A4;
        15'h1032: data = 12'h490;
        15'h1033: data = 12'h478;
        15'h1034: data = 12'h460;
        15'h1035: data = 12'h44D;
        15'h1036: data = 12'h432;
        15'h1037: data = 12'h419;
        15'h1038: data = 12'h401;
        15'h1039: data = 12'h3E8;
        15'h103A: data = 12'h3D4;
        15'h103B: data = 12'h3C5;
        15'h103C: data = 12'h3AA;
        15'h103D: data = 12'h38F;
        15'h103E: data = 12'h37F;
        15'h103F: data = 12'h363;
        15'h1040: data = 12'h351;
        15'h1041: data = 12'h337;
        15'h1042: data = 12'h324;
        15'h1043: data = 12'h30F;
        15'h1044: data = 12'h2F6;
        15'h1045: data = 12'h2E2;
        15'h1046: data = 12'h2CE;
        15'h1047: data = 12'h2B6;
        15'h1048: data = 12'h29E;
        15'h1049: data = 12'h285;
        15'h104A: data = 12'h275;
        15'h104B: data = 12'h25E;
        15'h104C: data = 12'h247;
        15'h104D: data = 12'h230;
        15'h104E: data = 12'h217;
        15'h104F: data = 12'h201;
        15'h1050: data = 12'h1ED;
        15'h1051: data = 12'h1D2;
        15'h1052: data = 12'h1BC;
        15'h1053: data = 12'h1A4;
        15'h1054: data = 12'h18E;
        15'h1055: data = 12'h178;
        15'h1056: data = 12'h161;
        15'h1057: data = 12'h14B;
        15'h1058: data = 12'h132;
        15'h1059: data = 12'h11C;
        15'h105A: data = 12'h105;
        15'h105B: data = 12'h0EE;
        15'h105C: data = 12'h0DA;
        15'h105D: data = 12'h0BC;
        15'h105E: data = 12'h0A6;
        15'h105F: data = 12'h090;
        15'h1060: data = 12'h07F;
        15'h1061: data = 12'h063;
        15'h1062: data = 12'h049;
        15'h1063: data = 12'h334;
        15'h1064: data = 12'h7CA;
        15'h1065: data = 12'h7B7;
        15'h1066: data = 12'h79F;
        15'h1067: data = 12'h78B;
        15'h1068: data = 12'h775;
        15'h1069: data = 12'h75F;
        15'h106A: data = 12'h749;
        15'h106B: data = 12'h735;
        15'h106C: data = 12'h71B;
        15'h106D: data = 12'h704;
        15'h106E: data = 12'h6EF;
        15'h106F: data = 12'h6DB;
        15'h1070: data = 12'h6C7;
        15'h1071: data = 12'h6B0;
        15'h1072: data = 12'h69A;
        15'h1073: data = 12'h688;
        15'h1074: data = 12'h66D;
        15'h1075: data = 12'h659;
        15'h1076: data = 12'h63E;
        15'h1077: data = 12'h631;
        15'h1078: data = 12'h617;
        15'h1079: data = 12'h601;
        15'h107A: data = 12'h5EB;
        15'h107B: data = 12'h5D4;
        15'h107C: data = 12'h5C2;
        15'h107D: data = 12'h5A8;
        15'h107E: data = 12'h594;
        15'h107F: data = 12'h57C;
        15'h1080: data = 12'h569;
        15'h1081: data = 12'h555;
        15'h1082: data = 12'h541;
        15'h1083: data = 12'h524;
        15'h1084: data = 12'h515;
        15'h1085: data = 12'h4F9;
        15'h1086: data = 12'h4E3;
        15'h1087: data = 12'h4D0;
        15'h1088: data = 12'h4BA;
        15'h1089: data = 12'h4A7;
        15'h108A: data = 12'h48D;
        15'h108B: data = 12'h47E;
        15'h108C: data = 12'h468;
        15'h108D: data = 12'h453;
        15'h108E: data = 12'h442;
        15'h108F: data = 12'h434;
        15'h1090: data = 12'h420;
        15'h1091: data = 12'h413;
        15'h1092: data = 12'h3FE;
        15'h1093: data = 12'h3EF;
        15'h1094: data = 12'h3E1;
        15'h1095: data = 12'h3D2;
        15'h1096: data = 12'h3C2;
        15'h1097: data = 12'h3B0;
        15'h1098: data = 12'h3A1;
        15'h1099: data = 12'h394;
        15'h109A: data = 12'h37D;
        15'h109B: data = 12'h36B;
        15'h109C: data = 12'h359;
        15'h109D: data = 12'h348;
        15'h109E: data = 12'h339;
        15'h109F: data = 12'h324;
        15'h10A0: data = 12'h311;
        15'h10A1: data = 12'h2FD;
        15'h10A2: data = 12'h2EE;
        15'h10A3: data = 12'h2DE;
        15'h10A4: data = 12'h2D1;
        15'h10A5: data = 12'h2C9;
        15'h10A6: data = 12'h2BB;
        15'h10A7: data = 12'h2AF;
        15'h10A8: data = 12'h2A4;
        15'h10A9: data = 12'h29C;
        15'h10AA: data = 12'h293;
        15'h10AB: data = 12'h284;
        15'h10AC: data = 12'h27C;
        15'h10AD: data = 12'h26E;
        15'h10AE: data = 12'h264;
        15'h10AF: data = 12'h256;
        15'h10B0: data = 12'h24B;
        15'h10B1: data = 12'h239;
        15'h10B2: data = 12'h22B;
        15'h10B3: data = 12'h21B;
        15'h10B4: data = 12'h210;
        15'h10B5: data = 12'h207;
        15'h10B6: data = 12'h1FD;
        15'h10B7: data = 12'h1EF;
        15'h10B8: data = 12'h1E8;
        15'h10B9: data = 12'h1E5;
        15'h10BA: data = 12'h1E0;
        15'h10BB: data = 12'h1DE;
        15'h10BC: data = 12'h1D8;
        15'h10BD: data = 12'h1CC;
        15'h10BE: data = 12'h1C8;
        15'h10BF: data = 12'h1C1;
        15'h10C0: data = 12'h1B9;
        15'h10C1: data = 12'h1AD;
        15'h10C2: data = 12'h1A1;
        15'h10C3: data = 12'h198;
        15'h10C4: data = 12'h192;
        15'h10C5: data = 12'h187;
        15'h10C6: data = 12'h182;
        15'h10C7: data = 12'h17F;
        15'h10C8: data = 12'h17F;
        15'h10C9: data = 12'h17A;
        15'h10CA: data = 12'h180;
        15'h10CB: data = 12'h17E;
        15'h10CC: data = 12'h17E;
        15'h10CD: data = 12'h176;
        15'h10CE: data = 12'h178;
        15'h10CF: data = 12'h175;
        15'h10D0: data = 12'h16B;
        15'h10D1: data = 12'h168;
        15'h10D2: data = 12'h161;
        15'h10D3: data = 12'h15F;
        15'h10D4: data = 12'h153;
        15'h10D5: data = 12'h156;
        15'h10D6: data = 12'h155;
        15'h10D7: data = 12'h154;
        15'h10D8: data = 12'h156;
        15'h10D9: data = 12'h15D;
        15'h10DA: data = 12'h161;
        15'h10DB: data = 12'h168;
        15'h10DC: data = 12'h16D;
        15'h10DD: data = 12'h16F;
        15'h10DE: data = 12'h16C;
        15'h10DF: data = 12'h16C;
        15'h10E0: data = 12'h173;
        15'h10E1: data = 12'h16D;
        15'h10E2: data = 12'h16D;
        15'h10E3: data = 12'h174;
        15'h10E4: data = 12'h16F;
        15'h10E5: data = 12'h177;
        15'h10E6: data = 12'h178;
        15'h10E7: data = 12'h17E;
        15'h10E8: data = 12'h188;
        15'h10E9: data = 12'h188;
        15'h10EA: data = 12'h194;
        15'h10EB: data = 12'h1A1;
        15'h10EC: data = 12'h1AB;
        15'h10ED: data = 12'h1B4;
        15'h10EE: data = 12'h1B2;
        15'h10EF: data = 12'h1BB;
        15'h10F0: data = 12'h1C3;
        15'h10F1: data = 12'h1C5;
        15'h10F2: data = 12'h1CA;
        15'h10F3: data = 12'h1CD;
        15'h10F4: data = 12'h1D2;
        15'h10F5: data = 12'h1D6;
        15'h10F6: data = 12'h1E0;
        15'h10F7: data = 12'h1E7;
        15'h10F8: data = 12'h1F6;
        15'h10F9: data = 12'h1FF;
        15'h10FA: data = 12'h20A;
        15'h10FB: data = 12'h213;
        15'h10FC: data = 12'h227;
        15'h10FD: data = 12'h234;
        15'h10FE: data = 12'h243;
        15'h10FF: data = 12'h24E;
        15'h1100: data = 12'h25F;
        15'h1101: data = 12'h264;
        15'h1102: data = 12'h272;
        15'h1103: data = 12'h275;
        15'h1104: data = 12'h283;
        15'h1105: data = 12'h28A;
        15'h1106: data = 12'h295;
        15'h1107: data = 12'h29E;
        15'h1108: data = 12'h2AE;
        15'h1109: data = 12'h2BD;
        15'h110A: data = 12'h2CA;
        15'h110B: data = 12'h2D6;
        15'h110C: data = 12'h2E6;
        15'h110D: data = 12'h2FC;
        15'h110E: data = 12'h30E;
        15'h110F: data = 12'h321;
        15'h1110: data = 12'h335;
        15'h1111: data = 12'h342;
        15'h1112: data = 12'h352;
        15'h1113: data = 12'h363;
        15'h1114: data = 12'h375;
        15'h1115: data = 12'h381;
        15'h1116: data = 12'h396;
        15'h1117: data = 12'h39E;
        15'h1118: data = 12'h3B4;
        15'h1119: data = 12'h3BF;
        15'h111A: data = 12'h3CC;
        15'h111B: data = 12'h3DF;
        15'h111C: data = 12'h3ED;
        15'h111D: data = 12'h3FC;
        15'h111E: data = 12'h412;
        15'h111F: data = 12'h423;
        15'h1120: data = 12'h435;
        15'h1121: data = 12'h44E;
        15'h1122: data = 12'h461;
        15'h1123: data = 12'h479;
        15'h1124: data = 12'h488;
        15'h1125: data = 12'h4A6;
        15'h1126: data = 12'h4B8;
        15'h1127: data = 12'h4D1;
        15'h1128: data = 12'h4E1;
        15'h1129: data = 12'h4F5;
        15'h112A: data = 12'h50A;
        15'h112B: data = 12'h51D;
        15'h112C: data = 12'h534;
        15'h112D: data = 12'h547;
        15'h112E: data = 12'h55A;
        15'h112F: data = 12'h568;
        15'h1130: data = 12'h576;
        15'h1131: data = 12'h58B;
        15'h1132: data = 12'h59D;
        15'h1133: data = 12'h5B1;
        15'h1134: data = 12'h5C8;
        15'h1135: data = 12'h5DF;
        15'h1136: data = 12'h5F5;
        15'h1137: data = 12'h60F;
        15'h1138: data = 12'h621;
        15'h1139: data = 12'h63B;
        15'h113A: data = 12'h65A;
        15'h113B: data = 12'h66D;
        15'h113C: data = 12'h68A;
        15'h113D: data = 12'h69C;
        15'h113E: data = 12'h6B8;
        15'h113F: data = 12'h6CC;
        15'h1140: data = 12'h6E3;
        15'h1141: data = 12'h6F9;
        15'h1142: data = 12'h711;
        15'h1143: data = 12'h726;
        15'h1144: data = 12'h73D;
        15'h1145: data = 12'h74E;
        15'h1146: data = 12'h762;
        15'h1147: data = 12'h775;
        15'h1148: data = 12'h78E;
        15'h1149: data = 12'h7A1;
        15'h114A: data = 12'h7B5;
        15'h114B: data = 12'h7CE;
        15'h114C: data = 12'h7E4;
        15'h114D: data = 12'h7FA;
        15'h114E: data = 12'h067;
        15'h114F: data = 12'h07E;
        15'h1150: data = 12'h095;
        15'h1151: data = 12'h0AA;
        15'h1152: data = 12'h0C3;
        15'h1153: data = 12'h0E4;
        15'h1154: data = 12'h0FD;
        15'h1155: data = 12'h110;
        15'h1156: data = 12'h127;
        15'h1157: data = 12'h144;
        15'h1158: data = 12'h157;
        15'h1159: data = 12'h16D;
        15'h115A: data = 12'h184;
        15'h115B: data = 12'h19C;
        15'h115C: data = 12'h1B9;
        15'h115D: data = 12'h1C7;
        15'h115E: data = 12'h1DE;
        15'h115F: data = 12'h1F7;
        15'h1160: data = 12'h20A;
        15'h1161: data = 12'h219;
        15'h1162: data = 12'h234;
        15'h1163: data = 12'h24B;
        15'h1164: data = 12'h262;
        15'h1165: data = 12'h275;
        15'h1166: data = 12'h285;
        15'h1167: data = 12'h2A3;
        15'h1168: data = 12'h2BA;
        15'h1169: data = 12'h2C7;
        15'h116A: data = 12'h2E9;
        15'h116B: data = 12'h2FB;
        15'h116C: data = 12'h31A;
        15'h116D: data = 12'h329;
        15'h116E: data = 12'h342;
        15'h116F: data = 12'h35B;
        15'h1170: data = 12'h373;
        15'h1171: data = 12'h38F;
        15'h1172: data = 12'h3A3;
        15'h1173: data = 12'h3BF;
        15'h1174: data = 12'h3D7;
        15'h1175: data = 12'h3EE;
        15'h1176: data = 12'h401;
        15'h1177: data = 12'h419;
        15'h1178: data = 12'h42F;
        15'h1179: data = 12'h445;
        15'h117A: data = 12'h458;
        15'h117B: data = 12'h46B;
        15'h117C: data = 12'h482;
        15'h117D: data = 12'h496;
        15'h117E: data = 12'h4AA;
        15'h117F: data = 12'h4BD;
        15'h1180: data = 12'h4CC;
        15'h1181: data = 12'h4E1;
        15'h1182: data = 12'h4F6;
        15'h1183: data = 12'h508;
        15'h1184: data = 12'h516;
        15'h1185: data = 12'h529;
        15'h1186: data = 12'h53E;
        15'h1187: data = 12'h54B;
        15'h1188: data = 12'h55F;
        15'h1189: data = 12'h56F;
        15'h118A: data = 12'h582;
        15'h118B: data = 12'h593;
        15'h118C: data = 12'h5A4;
        15'h118D: data = 12'h5BA;
        15'h118E: data = 12'h5C6;
        15'h118F: data = 12'h5D6;
        15'h1190: data = 12'h5E7;
        15'h1191: data = 12'h5FB;
        15'h1192: data = 12'h609;
        15'h1193: data = 12'h615;
        15'h1194: data = 12'h627;
        15'h1195: data = 12'h633;
        15'h1196: data = 12'h649;
        15'h1197: data = 12'h65D;
        15'h1198: data = 12'h66B;
        15'h1199: data = 12'h677;
        15'h119A: data = 12'h68F;
        15'h119B: data = 12'h69A;
        15'h119C: data = 12'h6A7;
        15'h119D: data = 12'h6B7;
        15'h119E: data = 12'h6C8;
        15'h119F: data = 12'h6D3;
        15'h11A0: data = 12'h6E3;
        15'h11A1: data = 12'h6F5;
        15'h11A2: data = 12'h6FD;
        15'h11A3: data = 12'h710;
        15'h11A4: data = 12'h720;
        15'h11A5: data = 12'h72C;
        15'h11A6: data = 12'h733;
        15'h11A7: data = 12'h73F;
        15'h11A8: data = 12'h74C;
        15'h11A9: data = 12'h75A;
        15'h11AA: data = 12'h768;
        15'h11AB: data = 12'h777;
        15'h11AC: data = 12'h77E;
        15'h11AD: data = 12'h78B;
        15'h11AE: data = 12'h792;
        15'h11AF: data = 12'h79B;
        15'h11B0: data = 12'h7A6;
        15'h11B1: data = 12'h7AD;
        15'h11B2: data = 12'h7BA;
        15'h11B3: data = 12'h7C3;
        15'h11B4: data = 12'h7CC;
        15'h11B5: data = 12'h7D0;
        15'h11B6: data = 12'h7D9;
        15'h11B7: data = 12'h7DE;
        15'h11B8: data = 12'h7E7;
        15'h11B9: data = 12'h7EE;
        15'h11BA: data = 12'h7F6;
        15'h11BB: data = 12'h7FA;
        15'h11BC: data = 12'h805;
        15'h11BD: data = 12'h805;
        15'h11BE: data = 12'h80A;
        15'h11BF: data = 12'h811;
        15'h11C0: data = 12'h894;
        15'h11C1: data = 12'h08F;
        15'h11C2: data = 12'h097;
        15'h11C3: data = 12'h09F;
        15'h11C4: data = 12'h09F;
        15'h11C5: data = 12'h0A7;
        15'h11C6: data = 12'h0A6;
        15'h11C7: data = 12'h0AD;
        15'h11C8: data = 12'h0AF;
        15'h11C9: data = 12'h0AE;
        15'h11CA: data = 12'h0B5;
        15'h11CB: data = 12'h0B7;
        15'h11CC: data = 12'h0B6;
        15'h11CD: data = 12'h0B6;
        15'h11CE: data = 12'h0BE;
        15'h11CF: data = 12'h0C2;
        15'h11D0: data = 12'h0C7;
        15'h11D1: data = 12'h0C4;
        15'h11D2: data = 12'h0C8;
        15'h11D3: data = 12'h0CB;
        15'h11D4: data = 12'h0D0;
        15'h11D5: data = 12'h0C9;
        15'h11D6: data = 12'h0CC;
        15'h11D7: data = 12'h0CF;
        15'h11D8: data = 12'h0CA;
        15'h11D9: data = 12'h0CA;
        15'h11DA: data = 12'h0C1;
        15'h11DB: data = 12'h0C0;
        15'h11DC: data = 12'h0B2;
        15'h11DD: data = 12'h0AE;
        15'h11DE: data = 12'h0A7;
        15'h11DF: data = 12'h0A3;
        15'h11E0: data = 12'h0A3;
        15'h11E1: data = 12'h0A6;
        15'h11E2: data = 12'h0A5;
        15'h11E3: data = 12'h0A0;
        15'h11E4: data = 12'h0A3;
        15'h11E5: data = 12'h09D;
        15'h11E6: data = 12'h096;
        15'h11E7: data = 12'h08A;
        15'h11E8: data = 12'h07F;
        15'h11E9: data = 12'h075;
        15'h11EA: data = 12'h06B;
        15'h11EB: data = 12'h064;
        15'h11EC: data = 12'h062;
        15'h11ED: data = 12'h05D;
        15'h11EE: data = 12'h060;
        15'h11EF: data = 12'h057;
        15'h11F0: data = 12'h04E;
        15'h11F1: data = 12'h040;
        15'h11F2: data = 12'h7C4;
        15'h11F3: data = 12'h7B0;
        15'h11F4: data = 12'h7A0;
        15'h11F5: data = 12'h792;
        15'h11F6: data = 12'h78A;
        15'h11F7: data = 12'h788;
        15'h11F8: data = 12'h77A;
        15'h11F9: data = 12'h772;
        15'h11FA: data = 12'h764;
        15'h11FB: data = 12'h751;
        15'h11FC: data = 12'h73E;
        15'h11FD: data = 12'h72F;
        15'h11FE: data = 12'h720;
        15'h11FF: data = 12'h713;
        15'h1200: data = 12'h709;
        15'h1201: data = 12'h704;
        15'h1202: data = 12'h6F9;
        15'h1203: data = 12'h6EB;
        15'h1204: data = 12'h6E5;
        15'h1205: data = 12'h6D2;
        15'h1206: data = 12'h6BD;
        15'h1207: data = 12'h6AA;
        15'h1208: data = 12'h696;
        15'h1209: data = 12'h685;
        15'h120A: data = 12'h676;
        15'h120B: data = 12'h66B;
        15'h120C: data = 12'h662;
        15'h120D: data = 12'h655;
        15'h120E: data = 12'h648;
        15'h120F: data = 12'h635;
        15'h1210: data = 12'h62C;
        15'h1211: data = 12'h614;
        15'h1212: data = 12'h603;
        15'h1213: data = 12'h5ED;
        15'h1214: data = 12'h5D3;
        15'h1215: data = 12'h5BE;
        15'h1216: data = 12'h5B1;
        15'h1217: data = 12'h5A1;
        15'h1218: data = 12'h58A;
        15'h1219: data = 12'h57D;
        15'h121A: data = 12'h56C;
        15'h121B: data = 12'h55D;
        15'h121C: data = 12'h554;
        15'h121D: data = 12'h541;
        15'h121E: data = 12'h52C;
        15'h121F: data = 12'h51C;
        15'h1220: data = 12'h508;
        15'h1221: data = 12'h4F5;
        15'h1222: data = 12'h4DD;
        15'h1223: data = 12'h4C9;
        15'h1224: data = 12'h4B6;
        15'h1225: data = 12'h49D;
        15'h1226: data = 12'h485;
        15'h1227: data = 12'h472;
        15'h1228: data = 12'h458;
        15'h1229: data = 12'h441;
        15'h122A: data = 12'h42D;
        15'h122B: data = 12'h415;
        15'h122C: data = 12'h3FD;
        15'h122D: data = 12'h3E6;
        15'h122E: data = 12'h3D3;
        15'h122F: data = 12'h3C0;
        15'h1230: data = 12'h3AC;
        15'h1231: data = 12'h390;
        15'h1232: data = 12'h37E;
        15'h1233: data = 12'h366;
        15'h1234: data = 12'h34F;
        15'h1235: data = 12'h33B;
        15'h1236: data = 12'h32B;
        15'h1237: data = 12'h315;
        15'h1238: data = 12'h2FB;
        15'h1239: data = 12'h2E9;
        15'h123A: data = 12'h2D8;
        15'h123B: data = 12'h2C1;
        15'h123C: data = 12'h2A6;
        15'h123D: data = 12'h28E;
        15'h123E: data = 12'h27A;
        15'h123F: data = 12'h265;
        15'h1240: data = 12'h24A;
        15'h1241: data = 12'h236;
        15'h1242: data = 12'h21C;
        15'h1243: data = 12'h205;
        15'h1244: data = 12'h1F2;
        15'h1245: data = 12'h1D8;
        15'h1246: data = 12'h1C0;
        15'h1247: data = 12'h1AA;
        15'h1248: data = 12'h195;
        15'h1249: data = 12'h17E;
        15'h124A: data = 12'h163;
        15'h124B: data = 12'h150;
        15'h124C: data = 12'h138;
        15'h124D: data = 12'h121;
        15'h124E: data = 12'h106;
        15'h124F: data = 12'h0F4;
        15'h1250: data = 12'h0DD;
        15'h1251: data = 12'h0C2;
        15'h1252: data = 12'h0A7;
        15'h1253: data = 12'h095;
        15'h1254: data = 12'h082;
        15'h1255: data = 12'h065;
        15'h1256: data = 12'h04D;
        15'h1257: data = 12'h47B;
        15'h1258: data = 12'h7CE;
        15'h1259: data = 12'h7BA;
        15'h125A: data = 12'h7A5;
        15'h125B: data = 12'h78E;
        15'h125C: data = 12'h776;
        15'h125D: data = 12'h761;
        15'h125E: data = 12'h74C;
        15'h125F: data = 12'h735;
        15'h1260: data = 12'h71E;
        15'h1261: data = 12'h709;
        15'h1262: data = 12'h6EF;
        15'h1263: data = 12'h6DD;
        15'h1264: data = 12'h6C7;
        15'h1265: data = 12'h6AE;
        15'h1266: data = 12'h698;
        15'h1267: data = 12'h687;
        15'h1268: data = 12'h669;
        15'h1269: data = 12'h659;
        15'h126A: data = 12'h63C;
        15'h126B: data = 12'h62C;
        15'h126C: data = 12'h614;
        15'h126D: data = 12'h5FA;
        15'h126E: data = 12'h5E5;
        15'h126F: data = 12'h5CE;
        15'h1270: data = 12'h5BF;
        15'h1271: data = 12'h5A2;
        15'h1272: data = 12'h58D;
        15'h1273: data = 12'h578;
        15'h1274: data = 12'h561;
        15'h1275: data = 12'h550;
        15'h1276: data = 12'h536;
        15'h1277: data = 12'h51F;
        15'h1278: data = 12'h50D;
        15'h1279: data = 12'h4F3;
        15'h127A: data = 12'h4DC;
        15'h127B: data = 12'h4CB;
        15'h127C: data = 12'h4B4;
        15'h127D: data = 12'h4A6;
        15'h127E: data = 12'h491;
        15'h127F: data = 12'h47F;
        15'h1280: data = 12'h46A;
        15'h1281: data = 12'h452;
        15'h1282: data = 12'h448;
        15'h1283: data = 12'h43B;
        15'h1284: data = 12'h427;
        15'h1285: data = 12'h417;
        15'h1286: data = 12'h401;
        15'h1287: data = 12'h3F7;
        15'h1288: data = 12'h3E9;
        15'h1289: data = 12'h3D4;
        15'h128A: data = 12'h3C2;
        15'h128B: data = 12'h3B4;
        15'h128C: data = 12'h39D;
        15'h128D: data = 12'h391;
        15'h128E: data = 12'h37C;
        15'h128F: data = 12'h36A;
        15'h1290: data = 12'h356;
        15'h1291: data = 12'h342;
        15'h1292: data = 12'h335;
        15'h1293: data = 12'h320;
        15'h1294: data = 12'h30D;
        15'h1295: data = 12'h2FF;
        15'h1296: data = 12'h2EF;
        15'h1297: data = 12'h2DF;
        15'h1298: data = 12'h2D1;
        15'h1299: data = 12'h2CC;
        15'h129A: data = 12'h2C2;
        15'h129B: data = 12'h2B4;
        15'h129C: data = 12'h2A7;
        15'h129D: data = 12'h2A1;
        15'h129E: data = 12'h291;
        15'h129F: data = 12'h285;
        15'h12A0: data = 12'h27F;
        15'h12A1: data = 12'h26C;
        15'h12A2: data = 12'h263;
        15'h12A3: data = 12'h24E;
        15'h12A4: data = 12'h243;
        15'h12A5: data = 12'h232;
        15'h12A6: data = 12'h225;
        15'h12A7: data = 12'h215;
        15'h12A8: data = 12'h20F;
        15'h12A9: data = 12'h20A;
        15'h12AA: data = 12'h200;
        15'h12AB: data = 12'h1F2;
        15'h12AC: data = 12'h1F1;
        15'h12AD: data = 12'h1EC;
        15'h12AE: data = 12'h1E8;
        15'h12AF: data = 12'h1E2;
        15'h12B0: data = 12'h1DC;
        15'h12B1: data = 12'h1CB;
        15'h12B2: data = 12'h1C6;
        15'h12B3: data = 12'h1BE;
        15'h12B4: data = 12'h1B4;
        15'h12B5: data = 12'h1A7;
        15'h12B6: data = 12'h19D;
        15'h12B7: data = 12'h194;
        15'h12B8: data = 12'h18C;
        15'h12B9: data = 12'h18A;
        15'h12BA: data = 12'h183;
        15'h12BB: data = 12'h186;
        15'h12BC: data = 12'h185;
        15'h12BD: data = 12'h180;
        15'h12BE: data = 12'h184;
        15'h12BF: data = 12'h180;
        15'h12C0: data = 12'h17F;
        15'h12C1: data = 12'h177;
        15'h12C2: data = 12'h178;
        15'h12C3: data = 12'h174;
        15'h12C4: data = 12'h166;
        15'h12C5: data = 12'h162;
        15'h12C6: data = 12'h15C;
        15'h12C7: data = 12'h15E;
        15'h12C8: data = 12'h152;
        15'h12C9: data = 12'h156;
        15'h12CA: data = 12'h158;
        15'h12CB: data = 12'h15B;
        15'h12CC: data = 12'h15F;
        15'h12CD: data = 12'h166;
        15'h12CE: data = 12'h168;
        15'h12CF: data = 12'h171;
        15'h12D0: data = 12'h16E;
        15'h12D1: data = 12'h16F;
        15'h12D2: data = 12'h16C;
        15'h12D3: data = 12'h16A;
        15'h12D4: data = 12'h16E;
        15'h12D5: data = 12'h168;
        15'h12D6: data = 12'h165;
        15'h12D7: data = 12'h16C;
        15'h12D8: data = 12'h168;
        15'h12D9: data = 12'h175;
        15'h12DA: data = 12'h17D;
        15'h12DB: data = 12'h185;
        15'h12DC: data = 12'h18C;
        15'h12DD: data = 12'h18F;
        15'h12DE: data = 12'h19A;
        15'h12DF: data = 12'h1A6;
        15'h12E0: data = 12'h1AC;
        15'h12E1: data = 12'h1B5;
        15'h12E2: data = 12'h1B1;
        15'h12E3: data = 12'h1B6;
        15'h12E4: data = 12'h1BE;
        15'h12E5: data = 12'h1C3;
        15'h12E6: data = 12'h1C7;
        15'h12E7: data = 12'h1CC;
        15'h12E8: data = 12'h1D2;
        15'h12E9: data = 12'h1D5;
        15'h12EA: data = 12'h1DF;
        15'h12EB: data = 12'h1EA;
        15'h12EC: data = 12'h1FA;
        15'h12ED: data = 12'h207;
        15'h12EE: data = 12'h214;
        15'h12EF: data = 12'h21C;
        15'h12F0: data = 12'h22D;
        15'h12F1: data = 12'h235;
        15'h12F2: data = 12'h247;
        15'h12F3: data = 12'h24E;
        15'h12F4: data = 12'h25C;
        15'h12F5: data = 12'h263;
        15'h12F6: data = 12'h270;
        15'h12F7: data = 12'h276;
        15'h12F8: data = 12'h27F;
        15'h12F9: data = 12'h284;
        15'h12FA: data = 12'h291;
        15'h12FB: data = 12'h29E;
        15'h12FC: data = 12'h2B2;
        15'h12FD: data = 12'h2BE;
        15'h12FE: data = 12'h2CA;
        15'h12FF: data = 12'h2DD;
        15'h1300: data = 12'h2EE;
        15'h1301: data = 12'h301;
        15'h1302: data = 12'h315;
        15'h1303: data = 12'h327;
        15'h1304: data = 12'h334;
        15'h1305: data = 12'h347;
        15'h1306: data = 12'h355;
        15'h1307: data = 12'h363;
        15'h1308: data = 12'h373;
        15'h1309: data = 12'h380;
        15'h130A: data = 12'h395;
        15'h130B: data = 12'h39B;
        15'h130C: data = 12'h3AF;
        15'h130D: data = 12'h3BB;
        15'h130E: data = 12'h3C9;
        15'h130F: data = 12'h3DC;
        15'h1310: data = 12'h3EA;
        15'h1311: data = 12'h3F8;
        15'h1312: data = 12'h416;
        15'h1313: data = 12'h429;
        15'h1314: data = 12'h43F;
        15'h1315: data = 12'h458;
        15'h1316: data = 12'h466;
        15'h1317: data = 12'h480;
        15'h1318: data = 12'h492;
        15'h1319: data = 12'h4AC;
        15'h131A: data = 12'h4BA;
        15'h131B: data = 12'h4D0;
        15'h131C: data = 12'h4E1;
        15'h131D: data = 12'h4F5;
        15'h131E: data = 12'h50C;
        15'h131F: data = 12'h518;
        15'h1320: data = 12'h52C;
        15'h1321: data = 12'h540;
        15'h1322: data = 12'h552;
        15'h1323: data = 12'h563;
        15'h1324: data = 12'h575;
        15'h1325: data = 12'h58C;
        15'h1326: data = 12'h59E;
        15'h1327: data = 12'h5B4;
        15'h1328: data = 12'h5CB;
        15'h1329: data = 12'h5E5;
        15'h132A: data = 12'h5FF;
        15'h132B: data = 12'h618;
        15'h132C: data = 12'h62C;
        15'h132D: data = 12'h646;
        15'h132E: data = 12'h65F;
        15'h132F: data = 12'h672;
        15'h1330: data = 12'h691;
        15'h1331: data = 12'h6A2;
        15'h1332: data = 12'h6B9;
        15'h1333: data = 12'h6CF;
        15'h1334: data = 12'h6E5;
        15'h1335: data = 12'h6F5;
        15'h1336: data = 12'h70D;
        15'h1337: data = 12'h722;
        15'h1338: data = 12'h736;
        15'h1339: data = 12'h747;
        15'h133A: data = 12'h75A;
        15'h133B: data = 12'h772;
        15'h133C: data = 12'h78D;
        15'h133D: data = 12'h7A1;
        15'h133E: data = 12'h7BB;
        15'h133F: data = 12'h7D2;
        15'h1340: data = 12'h7E7;
        15'h1341: data = 12'h802;
        15'h1342: data = 12'h071;
        15'h1343: data = 12'h08B;
        15'h1344: data = 12'h0A1;
        15'h1345: data = 12'h0B2;
        15'h1346: data = 12'h0D0;
        15'h1347: data = 12'h0E7;
        15'h1348: data = 12'h103;
        15'h1349: data = 12'h111;
        15'h134A: data = 12'h12C;
        15'h134B: data = 12'h142;
        15'h134C: data = 12'h156;
        15'h134D: data = 12'h16D;
        15'h134E: data = 12'h17F;
        15'h134F: data = 12'h195;
        15'h1350: data = 12'h1AF;
        15'h1351: data = 12'h1BF;
        15'h1352: data = 12'h1D5;
        15'h1353: data = 12'h1EB;
        15'h1354: data = 12'h205;
        15'h1355: data = 12'h212;
        15'h1356: data = 12'h22F;
        15'h1357: data = 12'h248;
        15'h1358: data = 12'h260;
        15'h1359: data = 12'h273;
        15'h135A: data = 12'h287;
        15'h135B: data = 12'h2A3;
        15'h135C: data = 12'h2BE;
        15'h135D: data = 12'h2D3;
        15'h135E: data = 12'h2EB;
        15'h135F: data = 12'h303;
        15'h1360: data = 12'h321;
        15'h1361: data = 12'h334;
        15'h1362: data = 12'h34B;
        15'h1363: data = 12'h368;
        15'h1364: data = 12'h37C;
        15'h1365: data = 12'h394;
        15'h1366: data = 12'h3A8;
        15'h1367: data = 12'h3C5;
        15'h1368: data = 12'h3D9;
        15'h1369: data = 12'h3EF;
        15'h136A: data = 12'h400;
        15'h136B: data = 12'h419;
        15'h136C: data = 12'h42D;
        15'h136D: data = 12'h445;
        15'h136E: data = 12'h454;
        15'h136F: data = 12'h469;
        15'h1370: data = 12'h47F;
        15'h1371: data = 12'h491;
        15'h1372: data = 12'h4AA;
        15'h1373: data = 12'h4BB;
        15'h1374: data = 12'h4C6;
        15'h1375: data = 12'h4DB;
        15'h1376: data = 12'h4F5;
        15'h1377: data = 12'h502;
        15'h1378: data = 12'h511;
        15'h1379: data = 12'h525;
        15'h137A: data = 12'h53C;
        15'h137B: data = 12'h546;
        15'h137C: data = 12'h55E;
        15'h137D: data = 12'h56A;
        15'h137E: data = 12'h57E;
        15'h137F: data = 12'h594;
        15'h1380: data = 12'h59E;
        15'h1381: data = 12'h5BB;
        15'h1382: data = 12'h5C4;
        15'h1383: data = 12'h5D6;
        15'h1384: data = 12'h5E9;
        15'h1385: data = 12'h5FB;
        15'h1386: data = 12'h60A;
        15'h1387: data = 12'h61A;
        15'h1388: data = 12'h62A;
        15'h1389: data = 12'h639;
        15'h138A: data = 12'h64F;
        15'h138B: data = 12'h65F;
        15'h138C: data = 12'h670;
        15'h138D: data = 12'h67F;
        15'h138E: data = 12'h694;
        15'h138F: data = 12'h69F;
        15'h1390: data = 12'h6B1;
        15'h1391: data = 12'h6BF;
        15'h1392: data = 12'h6CD;
        15'h1393: data = 12'h6DA;
        15'h1394: data = 12'h6E8;
        15'h1395: data = 12'h6F9;
        15'h1396: data = 12'h704;
        15'h1397: data = 12'h714;
        15'h1398: data = 12'h723;
        15'h1399: data = 12'h732;
        15'h139A: data = 12'h735;
        15'h139B: data = 12'h742;
        15'h139C: data = 12'h751;
        15'h139D: data = 12'h75D;
        15'h139E: data = 12'h767;
        15'h139F: data = 12'h777;
        15'h13A0: data = 12'h77F;
        15'h13A1: data = 12'h78B;
        15'h13A2: data = 12'h795;
        15'h13A3: data = 12'h79A;
        15'h13A4: data = 12'h7A3;
        15'h13A5: data = 12'h7AC;
        15'h13A6: data = 12'h7B8;
        15'h13A7: data = 12'h7C0;
        15'h13A8: data = 12'h7C5;
        15'h13A9: data = 12'h7CE;
        15'h13AA: data = 12'h7D3;
        15'h13AB: data = 12'h7DA;
        15'h13AC: data = 12'h7E4;
        15'h13AD: data = 12'h7E9;
        15'h13AE: data = 12'h7F3;
        15'h13AF: data = 12'h7FA;
        15'h13B0: data = 12'h7FF;
        15'h13B1: data = 12'h7FF;
        15'h13B2: data = 12'h805;
        15'h13B3: data = 12'h80A;
        15'h13B4: data = 12'h83D;
        15'h13B5: data = 12'h08A;
        15'h13B6: data = 12'h094;
        15'h13B7: data = 12'h099;
        15'h13B8: data = 12'h098;
        15'h13B9: data = 12'h09F;
        15'h13BA: data = 12'h09F;
        15'h13BB: data = 12'h0A9;
        15'h13BC: data = 12'h0A9;
        15'h13BD: data = 12'h0AA;
        15'h13BE: data = 12'h0B6;
        15'h13BF: data = 12'h0B6;
        15'h13C0: data = 12'h0B9;
        15'h13C1: data = 12'h0BB;
        15'h13C2: data = 12'h0C5;
        15'h13C3: data = 12'h0C4;
        15'h13C4: data = 12'h0C6;
        15'h13C5: data = 12'h0CD;
        15'h13C6: data = 12'h0D1;
        15'h13C7: data = 12'h0D3;
        15'h13C8: data = 12'h0D5;
        15'h13C9: data = 12'h0CD;
        15'h13CA: data = 12'h0CF;
        15'h13CB: data = 12'h0CD;
        15'h13CC: data = 12'h0C9;
        15'h13CD: data = 12'h0C5;
        15'h13CE: data = 12'h0BB;
        15'h13CF: data = 12'h0B5;
        15'h13D0: data = 12'h0AB;
        15'h13D1: data = 12'h0AB;
        15'h13D2: data = 12'h0A6;
        15'h13D3: data = 12'h0A6;
        15'h13D4: data = 12'h0A8;
        15'h13D5: data = 12'h0AE;
        15'h13D6: data = 12'h0B0;
        15'h13D7: data = 12'h0A7;
        15'h13D8: data = 12'h0A7;
        15'h13D9: data = 12'h09A;
        15'h13DA: data = 12'h092;
        15'h13DB: data = 12'h084;
        15'h13DC: data = 12'h075;
        15'h13DD: data = 12'h071;
        15'h13DE: data = 12'h06B;
        15'h13DF: data = 12'h06A;
        15'h13E0: data = 12'h068;
        15'h13E1: data = 12'h065;
        15'h13E2: data = 12'h05E;
        15'h13E3: data = 12'h058;
        15'h13E4: data = 12'h04B;
        15'h13E5: data = 12'h7C4;
        15'h13E6: data = 12'h7B2;
        15'h13E7: data = 12'h7AB;
        15'h13E8: data = 12'h79E;
        15'h13E9: data = 12'h796;
        15'h13EA: data = 12'h791;
        15'h13EB: data = 12'h78B;
        15'h13EC: data = 12'h77D;
        15'h13ED: data = 12'h76F;
        15'h13EE: data = 12'h75C;
        15'h13EF: data = 12'h74A;
        15'h13F0: data = 12'h736;
        15'h13F1: data = 12'h72F;
        15'h13F2: data = 12'h722;
        15'h13F3: data = 12'h718;
        15'h13F4: data = 12'h710;
        15'h13F5: data = 12'h708;
        15'h13F6: data = 12'h6FC;
        15'h13F7: data = 12'h6EC;
        15'h13F8: data = 12'h6E1;
        15'h13F9: data = 12'h6CC;
        15'h13FA: data = 12'h6B9;
        15'h13FB: data = 12'h6A8;
        15'h13FC: data = 12'h693;
        15'h13FD: data = 12'h684;
        15'h13FE: data = 12'h673;
        15'h13FF: data = 12'h669;
        15'h1400: data = 12'h661;
        15'h1401: data = 12'h655;
        15'h1402: data = 12'h645;
        15'h1403: data = 12'h638;
        15'h1404: data = 12'h62D;
        15'h1405: data = 12'h613;
        15'h1406: data = 12'h5FF;
        15'h1407: data = 12'h5EA;
        15'h1408: data = 12'h5D0;
        15'h1409: data = 12'h5BF;
        15'h140A: data = 12'h5B1;
        15'h140B: data = 12'h59F;
        15'h140C: data = 12'h58C;
        15'h140D: data = 12'h57F;
        15'h140E: data = 12'h56C;
        15'h140F: data = 12'h55F;
        15'h1410: data = 12'h552;
        15'h1411: data = 12'h541;
        15'h1412: data = 12'h52B;
        15'h1413: data = 12'h51D;
        15'h1414: data = 12'h50A;
        15'h1415: data = 12'h4F6;
        15'h1416: data = 12'h4DB;
        15'h1417: data = 12'h4CB;
        15'h1418: data = 12'h4B7;
        15'h1419: data = 12'h49D;
        15'h141A: data = 12'h487;
        15'h141B: data = 12'h472;
        15'h141C: data = 12'h458;
        15'h141D: data = 12'h443;
        15'h141E: data = 12'h42E;
        15'h141F: data = 12'h414;
        15'h1420: data = 12'h400;
        15'h1421: data = 12'h3E4;
        15'h1422: data = 12'h3D3;
        15'h1423: data = 12'h3C0;
        15'h1424: data = 12'h3A9;
        15'h1425: data = 12'h391;
        15'h1426: data = 12'h37C;
        15'h1427: data = 12'h363;
        15'h1428: data = 12'h34E;
        15'h1429: data = 12'h338;
        15'h142A: data = 12'h328;
        15'h142B: data = 12'h313;
        15'h142C: data = 12'h2FA;
        15'h142D: data = 12'h2E5;
        15'h142E: data = 12'h2D1;
        15'h142F: data = 12'h2BF;
        15'h1430: data = 12'h2A5;
        15'h1431: data = 12'h28C;
        15'h1432: data = 12'h27A;
        15'h1433: data = 12'h264;
        15'h1434: data = 12'h24A;
        15'h1435: data = 12'h232;
        15'h1436: data = 12'h21A;
        15'h1437: data = 12'h204;
        15'h1438: data = 12'h1F3;
        15'h1439: data = 12'h1D6;
        15'h143A: data = 12'h1BD;
        15'h143B: data = 12'h1A8;
        15'h143C: data = 12'h193;
        15'h143D: data = 12'h178;
        15'h143E: data = 12'h165;
        15'h143F: data = 12'h14C;
        15'h1440: data = 12'h134;
        15'h1441: data = 12'h11C;
        15'h1442: data = 12'h107;
        15'h1443: data = 12'h0F0;
        15'h1444: data = 12'h0DB;
        15'h1445: data = 12'h0C1;
        15'h1446: data = 12'h0A6;
        15'h1447: data = 12'h08F;
        15'h1448: data = 12'h081;
        15'h1449: data = 12'h065;
        15'h144A: data = 12'h04B;
        15'h144B: data = 12'h7E0;
        15'h144C: data = 12'h7CD;
        15'h144D: data = 12'h7B9;
        15'h144E: data = 12'h7A4;
        15'h144F: data = 12'h78E;
        15'h1450: data = 12'h777;
        15'h1451: data = 12'h75D;
        15'h1452: data = 12'h74B;
        15'h1453: data = 12'h737;
        15'h1454: data = 12'h720;
        15'h1455: data = 12'h70A;
        15'h1456: data = 12'h6EF;
        15'h1457: data = 12'h6D7;
        15'h1458: data = 12'h6C3;
        15'h1459: data = 12'h6AC;
        15'h145A: data = 12'h696;
        15'h145B: data = 12'h685;
        15'h145C: data = 12'h66B;
        15'h145D: data = 12'h657;
        15'h145E: data = 12'h63E;
        15'h145F: data = 12'h62C;
        15'h1460: data = 12'h615;
        15'h1461: data = 12'h5FD;
        15'h1462: data = 12'h5E6;
        15'h1463: data = 12'h5D3;
        15'h1464: data = 12'h5C1;
        15'h1465: data = 12'h5A5;
        15'h1466: data = 12'h58E;
        15'h1467: data = 12'h576;
        15'h1468: data = 12'h564;
        15'h1469: data = 12'h550;
        15'h146A: data = 12'h539;
        15'h146B: data = 12'h51D;
        15'h146C: data = 12'h50C;
        15'h146D: data = 12'h4F8;
        15'h146E: data = 12'h4DF;
        15'h146F: data = 12'h4D0;
        15'h1470: data = 12'h4B5;
        15'h1471: data = 12'h4A3;
        15'h1472: data = 12'h490;
        15'h1473: data = 12'h47E;
        15'h1474: data = 12'h469;
        15'h1475: data = 12'h454;
        15'h1476: data = 12'h445;
        15'h1477: data = 12'h438;
        15'h1478: data = 12'h423;
        15'h1479: data = 12'h416;
        15'h147A: data = 12'h400;
        15'h147B: data = 12'h3F2;
        15'h147C: data = 12'h3E8;
        15'h147D: data = 12'h3D2;
        15'h147E: data = 12'h3C1;
        15'h147F: data = 12'h3B3;
        15'h1480: data = 12'h3A1;
        15'h1481: data = 12'h394;
        15'h1482: data = 12'h380;
        15'h1483: data = 12'h36A;
        15'h1484: data = 12'h357;
        15'h1485: data = 12'h347;
        15'h1486: data = 12'h335;
        15'h1487: data = 12'h322;
        15'h1488: data = 12'h30C;
        15'h1489: data = 12'h2FB;
        15'h148A: data = 12'h2EF;
        15'h148B: data = 12'h2E1;
        15'h148C: data = 12'h2D0;
        15'h148D: data = 12'h2CB;
        15'h148E: data = 12'h2C0;
        15'h148F: data = 12'h2B2;
        15'h1490: data = 12'h2A8;
        15'h1491: data = 12'h2A0;
        15'h1492: data = 12'h294;
        15'h1493: data = 12'h285;
        15'h1494: data = 12'h27B;
        15'h1495: data = 12'h26F;
        15'h1496: data = 12'h265;
        15'h1497: data = 12'h253;
        15'h1498: data = 12'h243;
        15'h1499: data = 12'h234;
        15'h149A: data = 12'h228;
        15'h149B: data = 12'h216;
        15'h149C: data = 12'h20E;
        15'h149D: data = 12'h208;
        15'h149E: data = 12'h1FF;
        15'h149F: data = 12'h1F2;
        15'h14A0: data = 12'h1F0;
        15'h14A1: data = 12'h1EA;
        15'h14A2: data = 12'h1E3;
        15'h14A3: data = 12'h1E1;
        15'h14A4: data = 12'h1D7;
        15'h14A5: data = 12'h1CD;
        15'h14A6: data = 12'h1C6;
        15'h14A7: data = 12'h1C1;
        15'h14A8: data = 12'h1B7;
        15'h14A9: data = 12'h1AB;
        15'h14AA: data = 12'h19C;
        15'h14AB: data = 12'h197;
        15'h14AC: data = 12'h194;
        15'h14AD: data = 12'h188;
        15'h14AE: data = 12'h184;
        15'h14AF: data = 12'h183;
        15'h14B0: data = 12'h184;
        15'h14B1: data = 12'h17F;
        15'h14B2: data = 12'h184;
        15'h14B3: data = 12'h180;
        15'h14B4: data = 12'h17F;
        15'h14B5: data = 12'h179;
        15'h14B6: data = 12'h177;
        15'h14B7: data = 12'h175;
        15'h14B8: data = 12'h168;
        15'h14B9: data = 12'h164;
        15'h14BA: data = 12'h160;
        15'h14BB: data = 12'h15D;
        15'h14BC: data = 12'h152;
        15'h14BD: data = 12'h156;
        15'h14BE: data = 12'h157;
        15'h14BF: data = 12'h15C;
        15'h14C0: data = 12'h15C;
        15'h14C1: data = 12'h163;
        15'h14C2: data = 12'h164;
        15'h14C3: data = 12'h16C;
        15'h14C4: data = 12'h171;
        15'h14C5: data = 12'h16F;
        15'h14C6: data = 12'h170;
        15'h14C7: data = 12'h16B;
        15'h14C8: data = 12'h171;
        15'h14C9: data = 12'h16F;
        15'h14CA: data = 12'h169;
        15'h14CB: data = 12'h16C;
        15'h14CC: data = 12'h16C;
        15'h14CD: data = 12'h173;
        15'h14CE: data = 12'h17D;
        15'h14CF: data = 12'h17F;
        15'h14D0: data = 12'h18B;
        15'h14D1: data = 12'h18F;
        15'h14D2: data = 12'h19B;
        15'h14D3: data = 12'h1A1;
        15'h14D4: data = 12'h1AA;
        15'h14D5: data = 12'h1B5;
        15'h14D6: data = 12'h1B3;
        15'h14D7: data = 12'h1BB;
        15'h14D8: data = 12'h1C1;
        15'h14D9: data = 12'h1C6;
        15'h14DA: data = 12'h1CA;
        15'h14DB: data = 12'h1CC;
        15'h14DC: data = 12'h1D3;
        15'h14DD: data = 12'h1DA;
        15'h14DE: data = 12'h1DF;
        15'h14DF: data = 12'h1EB;
        15'h14E0: data = 12'h1F8;
        15'h14E1: data = 12'h202;
        15'h14E2: data = 12'h211;
        15'h14E3: data = 12'h21B;
        15'h14E4: data = 12'h22D;
        15'h14E5: data = 12'h236;
        15'h14E6: data = 12'h248;
        15'h14E7: data = 12'h24D;
        15'h14E8: data = 12'h25E;
        15'h14E9: data = 12'h266;
        15'h14EA: data = 12'h274;
        15'h14EB: data = 12'h27A;
        15'h14EC: data = 12'h283;
        15'h14ED: data = 12'h28A;
        15'h14EE: data = 12'h293;
        15'h14EF: data = 12'h2A1;
        15'h14F0: data = 12'h2AF;
        15'h14F1: data = 12'h2BF;
        15'h14F2: data = 12'h2CC;
        15'h14F3: data = 12'h2D9;
        15'h14F4: data = 12'h2EB;
        15'h14F5: data = 12'h2FD;
        15'h14F6: data = 12'h313;
        15'h14F7: data = 12'h323;
        15'h14F8: data = 12'h336;
        15'h14F9: data = 12'h345;
        15'h14FA: data = 12'h356;
        15'h14FB: data = 12'h364;
        15'h14FC: data = 12'h372;
        15'h14FD: data = 12'h380;
        15'h14FE: data = 12'h396;
        15'h14FF: data = 12'h39F;
        15'h1500: data = 12'h3B4;
        15'h1501: data = 12'h3BC;
        15'h1502: data = 12'h3CA;
        15'h1503: data = 12'h3DC;
        15'h1504: data = 12'h3EE;
        15'h1505: data = 12'h3FC;
        15'h1506: data = 12'h410;
        15'h1507: data = 12'h425;
        15'h1508: data = 12'h433;
        15'h1509: data = 12'h44F;
        15'h150A: data = 12'h464;
        15'h150B: data = 12'h47D;
        15'h150C: data = 12'h48C;
        15'h150D: data = 12'h4A5;
        15'h150E: data = 12'h4B9;
        15'h150F: data = 12'h4D2;
        15'h1510: data = 12'h4E0;
        15'h1511: data = 12'h4F3;
        15'h1512: data = 12'h50C;
        15'h1513: data = 12'h51C;
        15'h1514: data = 12'h52D;
        15'h1515: data = 12'h543;
        15'h1516: data = 12'h558;
        15'h1517: data = 12'h566;
        15'h1518: data = 12'h576;
        15'h1519: data = 12'h589;
        15'h151A: data = 12'h59E;
        15'h151B: data = 12'h5B5;
        15'h151C: data = 12'h5C8;
        15'h151D: data = 12'h5E0;
        15'h151E: data = 12'h5F9;
        15'h151F: data = 12'h613;
        15'h1520: data = 12'h625;
        15'h1521: data = 12'h640;
        15'h1522: data = 12'h65D;
        15'h1523: data = 12'h673;
        15'h1524: data = 12'h68F;
        15'h1525: data = 12'h6A1;
        15'h1526: data = 12'h6B7;
        15'h1527: data = 12'h6D3;
        15'h1528: data = 12'h6E2;
        15'h1529: data = 12'h6F8;
        15'h152A: data = 12'h70F;
        15'h152B: data = 12'h727;
        15'h152C: data = 12'h73B;
        15'h152D: data = 12'h74E;
        15'h152E: data = 12'h75F;
        15'h152F: data = 12'h775;
        15'h1530: data = 12'h78D;
        15'h1531: data = 12'h7A0;
        15'h1532: data = 12'h7B7;
        15'h1533: data = 12'h7CE;
        15'h1534: data = 12'h7E5;
        15'h1535: data = 12'h7FD;
        15'h1536: data = 12'h06A;
        15'h1537: data = 12'h085;
        15'h1538: data = 12'h09D;
        15'h1539: data = 12'h0AC;
        15'h153A: data = 12'h0CB;
        15'h153B: data = 12'h0E9;
        15'h153C: data = 12'h0FE;
        15'h153D: data = 12'h112;
        15'h153E: data = 12'h12C;
        15'h153F: data = 12'h143;
        15'h1540: data = 12'h159;
        15'h1541: data = 12'h170;
        15'h1542: data = 12'h182;
        15'h1543: data = 12'h19C;
        15'h1544: data = 12'h1B5;
        15'h1545: data = 12'h1C0;
        15'h1546: data = 12'h1DA;
        15'h1547: data = 12'h1F1;
        15'h1548: data = 12'h207;
        15'h1549: data = 12'h217;
        15'h154A: data = 12'h230;
        15'h154B: data = 12'h249;
        15'h154C: data = 12'h262;
        15'h154D: data = 12'h275;
        15'h154E: data = 12'h288;
        15'h154F: data = 12'h2A4;
        15'h1550: data = 12'h2BD;
        15'h1551: data = 12'h2CE;
        15'h1552: data = 12'h2EA;
        15'h1553: data = 12'h2FE;
        15'h1554: data = 12'h31B;
        15'h1555: data = 12'h32D;
        15'h1556: data = 12'h348;
        15'h1557: data = 12'h361;
        15'h1558: data = 12'h376;
        15'h1559: data = 12'h391;
        15'h155A: data = 12'h3A8;
        15'h155B: data = 12'h3C3;
        15'h155C: data = 12'h3D6;
        15'h155D: data = 12'h3EF;
        15'h155E: data = 12'h404;
        15'h155F: data = 12'h419;
        15'h1560: data = 12'h42F;
        15'h1561: data = 12'h449;
        15'h1562: data = 12'h456;
        15'h1563: data = 12'h46A;
        15'h1564: data = 12'h482;
        15'h1565: data = 12'h495;
        15'h1566: data = 12'h4A9;
        15'h1567: data = 12'h4BC;
        15'h1568: data = 12'h4CA;
        15'h1569: data = 12'h4E3;
        15'h156A: data = 12'h4F8;
        15'h156B: data = 12'h50F;
        15'h156C: data = 12'h514;
        15'h156D: data = 12'h528;
        15'h156E: data = 12'h540;
        15'h156F: data = 12'h549;
        15'h1570: data = 12'h564;
        15'h1571: data = 12'h570;
        15'h1572: data = 12'h585;
        15'h1573: data = 12'h594;
        15'h1574: data = 12'h5A3;
        15'h1575: data = 12'h5B9;
        15'h1576: data = 12'h5C5;
        15'h1577: data = 12'h5D5;
        15'h1578: data = 12'h5E7;
        15'h1579: data = 12'h5F8;
        15'h157A: data = 12'h60A;
        15'h157B: data = 12'h617;
        15'h157C: data = 12'h627;
        15'h157D: data = 12'h635;
        15'h157E: data = 12'h648;
        15'h157F: data = 12'h65C;
        15'h1580: data = 12'h66D;
        15'h1581: data = 12'h676;
        15'h1582: data = 12'h68D;
        15'h1583: data = 12'h69C;
        15'h1584: data = 12'h6A4;
        15'h1585: data = 12'h6B6;
        15'h1586: data = 12'h6C6;
        15'h1587: data = 12'h6D2;
        15'h1588: data = 12'h6E1;
        15'h1589: data = 12'h6F2;
        15'h158A: data = 12'h6FB;
        15'h158B: data = 12'h70C;
        15'h158C: data = 12'h71A;
        15'h158D: data = 12'h72D;
        15'h158E: data = 12'h732;
        15'h158F: data = 12'h73F;
        15'h1590: data = 12'h74D;
        15'h1591: data = 12'h75B;
        15'h1592: data = 12'h763;
        15'h1593: data = 12'h771;
        15'h1594: data = 12'h77D;
        15'h1595: data = 12'h78B;
        15'h1596: data = 12'h792;
        15'h1597: data = 12'h79D;
        15'h1598: data = 12'h7A3;
        15'h1599: data = 12'h7AF;
        15'h159A: data = 12'h7BA;
        15'h159B: data = 12'h7C1;
        15'h159C: data = 12'h7C9;
        15'h159D: data = 12'h7D0;
        15'h159E: data = 12'h7D9;
        15'h159F: data = 12'h7E0;
        15'h15A0: data = 12'h7E7;
        15'h15A1: data = 12'h7ED;
        15'h15A2: data = 12'h7F6;
        15'h15A3: data = 12'h7FE;
        15'h15A4: data = 12'h806;
        15'h15A5: data = 12'h806;
        15'h15A6: data = 12'h809;
        15'h15A7: data = 12'h813;
        15'h15A8: data = 12'h876;
        15'h15A9: data = 12'h090;
        15'h15AA: data = 12'h09C;
        15'h15AB: data = 12'h09F;
        15'h15AC: data = 12'h0A2;
        15'h15AD: data = 12'h0A9;
        15'h15AE: data = 12'h0A7;
        15'h15AF: data = 12'h0AE;
        15'h15B0: data = 12'h0B0;
        15'h15B1: data = 12'h0B2;
        15'h15B2: data = 12'h0B7;
        15'h15B3: data = 12'h0B8;
        15'h15B4: data = 12'h0B5;
        15'h15B5: data = 12'h0B5;
        15'h15B6: data = 12'h0BD;
        15'h15B7: data = 12'h0BE;
        15'h15B8: data = 12'h0C1;
        15'h15B9: data = 12'h0C4;
        15'h15BA: data = 12'h0C7;
        15'h15BB: data = 12'h0CA;
        15'h15BC: data = 12'h0D1;
        15'h15BD: data = 12'h0C9;
        15'h15BE: data = 12'h0CC;
        15'h15BF: data = 12'h0CE;
        15'h15C0: data = 12'h0CD;
        15'h15C1: data = 12'h0CF;
        15'h15C2: data = 12'h0C7;
        15'h15C3: data = 12'h0C6;
        15'h15C4: data = 12'h0B7;
        15'h15C5: data = 12'h0B5;
        15'h15C6: data = 12'h0A6;
        15'h15C7: data = 12'h0A4;
        15'h15C8: data = 12'h09F;
        15'h15C9: data = 12'h0A5;
        15'h15CA: data = 12'h0A3;
        15'h15CB: data = 12'h0A1;
        15'h15CC: data = 12'h0A5;
        15'h15CD: data = 12'h0A1;
        15'h15CE: data = 12'h098;
        15'h15CF: data = 12'h08D;
        15'h15D0: data = 12'h080;
        15'h15D1: data = 12'h07B;
        15'h15D2: data = 12'h06F;
        15'h15D3: data = 12'h066;
        15'h15D4: data = 12'h060;
        15'h15D5: data = 12'h05C;
        15'h15D6: data = 12'h05C;
        15'h15D7: data = 12'h058;
        15'h15D8: data = 12'h051;
        15'h15D9: data = 12'h1B9;
        15'h15DA: data = 12'h7C1;
        15'h15DB: data = 12'h7AF;
        15'h15DC: data = 12'h79F;
        15'h15DD: data = 12'h791;
        15'h15DE: data = 12'h786;
        15'h15DF: data = 12'h785;
        15'h15E0: data = 12'h779;
        15'h15E1: data = 12'h775;
        15'h15E2: data = 12'h766;
        15'h15E3: data = 12'h75A;
        15'h15E4: data = 12'h743;
        15'h15E5: data = 12'h733;
        15'h15E6: data = 12'h724;
        15'h15E7: data = 12'h715;
        15'h15E8: data = 12'h709;
        15'h15E9: data = 12'h703;
        15'h15EA: data = 12'h6FA;
        15'h15EB: data = 12'h6EC;
        15'h15EC: data = 12'h6E5;
        15'h15ED: data = 12'h6D4;
        15'h15EE: data = 12'h6C0;
        15'h15EF: data = 12'h6AD;
        15'h15F0: data = 12'h698;
        15'h15F1: data = 12'h688;
        15'h15F2: data = 12'h677;
        15'h15F3: data = 12'h668;
        15'h15F4: data = 12'h65A;
        15'h15F5: data = 12'h64F;
        15'h15F6: data = 12'h645;
        15'h15F7: data = 12'h639;
        15'h15F8: data = 12'h62C;
        15'h15F9: data = 12'h617;
        15'h15FA: data = 12'h604;
        15'h15FB: data = 12'h5F9;
        15'h15FC: data = 12'h5DB;
        15'h15FD: data = 12'h5C3;
        15'h15FE: data = 12'h5B4;
        15'h15FF: data = 12'h5A3;
        15'h1600: data = 12'h58A;
        15'h1601: data = 12'h57C;
        15'h1602: data = 12'h567;
        15'h1603: data = 12'h559;
        15'h1604: data = 12'h54E;
        15'h1605: data = 12'h540;
        15'h1606: data = 12'h52C;
        15'h1607: data = 12'h51D;
        15'h1608: data = 12'h50B;
        15'h1609: data = 12'h4F7;
        15'h160A: data = 12'h4DF;
        15'h160B: data = 12'h4CC;
        15'h160C: data = 12'h4B8;
        15'h160D: data = 12'h4A4;
        15'h160E: data = 12'h490;
        15'h160F: data = 12'h476;
        15'h1610: data = 12'h45B;
        15'h1611: data = 12'h449;
        15'h1612: data = 12'h431;
        15'h1613: data = 12'h416;
        15'h1614: data = 12'h3FF;
        15'h1615: data = 12'h3E9;
        15'h1616: data = 12'h3D3;
        15'h1617: data = 12'h3BF;
        15'h1618: data = 12'h3AA;
        15'h1619: data = 12'h392;
        15'h161A: data = 12'h37D;
        15'h161B: data = 12'h364;
        15'h161C: data = 12'h34E;
        15'h161D: data = 12'h339;
        15'h161E: data = 12'h326;
        15'h161F: data = 12'h314;
        15'h1620: data = 12'h2F7;
        15'h1621: data = 12'h2E7;
        15'h1622: data = 12'h2D0;
        15'h1623: data = 12'h2BC;
        15'h1624: data = 12'h2A5;
        15'h1625: data = 12'h28B;
        15'h1626: data = 12'h27C;
        15'h1627: data = 12'h263;
        15'h1628: data = 12'h248;
        15'h1629: data = 12'h237;
        15'h162A: data = 12'h21C;
        15'h162B: data = 12'h207;
        15'h162C: data = 12'h1F3;
        15'h162D: data = 12'h1D8;
        15'h162E: data = 12'h1BE;
        15'h162F: data = 12'h1AA;
        15'h1630: data = 12'h197;
        15'h1631: data = 12'h17D;
        15'h1632: data = 12'h164;
        15'h1633: data = 12'h14F;
        15'h1634: data = 12'h137;
        15'h1635: data = 12'h11E;
        15'h1636: data = 12'h108;
        15'h1637: data = 12'h0F3;
        15'h1638: data = 12'h0E0;
        15'h1639: data = 12'h0C1;
        15'h163A: data = 12'h0A6;
        15'h163B: data = 12'h093;
        15'h163C: data = 12'h080;
        15'h163D: data = 12'h067;
        15'h163E: data = 12'h04D;
        15'h163F: data = 12'h40D;
        15'h1640: data = 12'h7CE;
        15'h1641: data = 12'h7BB;
        15'h1642: data = 12'h7A5;
        15'h1643: data = 12'h790;
        15'h1644: data = 12'h778;
        15'h1645: data = 12'h75E;
        15'h1646: data = 12'h74E;
        15'h1647: data = 12'h735;
        15'h1648: data = 12'h71D;
        15'h1649: data = 12'h706;
        15'h164A: data = 12'h6EC;
        15'h164B: data = 12'h6D9;
        15'h164C: data = 12'h6C6;
        15'h164D: data = 12'h6B2;
        15'h164E: data = 12'h699;
        15'h164F: data = 12'h685;
        15'h1650: data = 12'h669;
        15'h1651: data = 12'h65A;
        15'h1652: data = 12'h63F;
        15'h1653: data = 12'h62D;
        15'h1654: data = 12'h616;
        15'h1655: data = 12'h5FE;
        15'h1656: data = 12'h5E9;
        15'h1657: data = 12'h5D2;
        15'h1658: data = 12'h5C0;
        15'h1659: data = 12'h5A6;
        15'h165A: data = 12'h590;
        15'h165B: data = 12'h579;
        15'h165C: data = 12'h568;
        15'h165D: data = 12'h552;
        15'h165E: data = 12'h53A;
        15'h165F: data = 12'h520;
        15'h1660: data = 12'h50D;
        15'h1661: data = 12'h4F6;
        15'h1662: data = 12'h4DC;
        15'h1663: data = 12'h4CC;
        15'h1664: data = 12'h4B8;
        15'h1665: data = 12'h4A7;
        15'h1666: data = 12'h490;
        15'h1667: data = 12'h47E;
        15'h1668: data = 12'h466;
        15'h1669: data = 12'h452;
        15'h166A: data = 12'h444;
        15'h166B: data = 12'h437;
        15'h166C: data = 12'h421;
        15'h166D: data = 12'h412;
        15'h166E: data = 12'h400;
        15'h166F: data = 12'h3F4;
        15'h1670: data = 12'h3E9;
        15'h1671: data = 12'h3D4;
        15'h1672: data = 12'h3C3;
        15'h1673: data = 12'h3B2;
        15'h1674: data = 12'h39F;
        15'h1675: data = 12'h392;
        15'h1676: data = 12'h37C;
        15'h1677: data = 12'h36C;
        15'h1678: data = 12'h35A;
        15'h1679: data = 12'h345;
        15'h167A: data = 12'h335;
        15'h167B: data = 12'h323;
        15'h167C: data = 12'h30E;
        15'h167D: data = 12'h2FC;
        15'h167E: data = 12'h2F0;
        15'h167F: data = 12'h2E1;
        15'h1680: data = 12'h2D2;
        15'h1681: data = 12'h2C9;
        15'h1682: data = 12'h2BE;
        15'h1683: data = 12'h2B1;
        15'h1684: data = 12'h2A7;
        15'h1685: data = 12'h29F;
        15'h1686: data = 12'h294;
        15'h1687: data = 12'h285;
        15'h1688: data = 12'h281;
        15'h1689: data = 12'h26D;
        15'h168A: data = 12'h263;
        15'h168B: data = 12'h253;
        15'h168C: data = 12'h248;
        15'h168D: data = 12'h233;
        15'h168E: data = 12'h229;
        15'h168F: data = 12'h218;
        15'h1690: data = 12'h20C;
        15'h1691: data = 12'h205;
        15'h1692: data = 12'h1FF;
        15'h1693: data = 12'h1EF;
        15'h1694: data = 12'h1EB;
        15'h1695: data = 12'h1EA;
        15'h1696: data = 12'h1E6;
        15'h1697: data = 12'h1E0;
        15'h1698: data = 12'h1D9;
        15'h1699: data = 12'h1CE;
        15'h169A: data = 12'h1C6;
        15'h169B: data = 12'h1C1;
        15'h169C: data = 12'h1B8;
        15'h169D: data = 12'h1AC;
        15'h169E: data = 12'h1A0;
        15'h169F: data = 12'h198;
        15'h16A0: data = 12'h195;
        15'h16A1: data = 12'h18A;
        15'h16A2: data = 12'h184;
        15'h16A3: data = 12'h185;
        15'h16A4: data = 12'h180;
        15'h16A5: data = 12'h17F;
        15'h16A6: data = 12'h183;
        15'h16A7: data = 12'h17D;
        15'h16A8: data = 12'h17D;
        15'h16A9: data = 12'h178;
        15'h16AA: data = 12'h176;
        15'h16AB: data = 12'h175;
        15'h16AC: data = 12'h16A;
        15'h16AD: data = 12'h168;
        15'h16AE: data = 12'h161;
        15'h16AF: data = 12'h15D;
        15'h16B0: data = 12'h155;
        15'h16B1: data = 12'h155;
        15'h16B2: data = 12'h153;
        15'h16B3: data = 12'h157;
        15'h16B4: data = 12'h15D;
        15'h16B5: data = 12'h160;
        15'h16B6: data = 12'h165;
        15'h16B7: data = 12'h16D;
        15'h16B8: data = 12'h16D;
        15'h16B9: data = 12'h16F;
        15'h16BA: data = 12'h16D;
        15'h16BB: data = 12'h16B;
        15'h16BC: data = 12'h170;
        15'h16BD: data = 12'h16D;
        15'h16BE: data = 12'h16B;
        15'h16BF: data = 12'h16F;
        15'h16C0: data = 12'h16E;
        15'h16C1: data = 12'h172;
        15'h16C2: data = 12'h179;
        15'h16C3: data = 12'h17B;
        15'h16C4: data = 12'h187;
        15'h16C5: data = 12'h18B;
        15'h16C6: data = 12'h198;
        15'h16C7: data = 12'h1A4;
        15'h16C8: data = 12'h1AB;
        15'h16C9: data = 12'h1B2;
        15'h16CA: data = 12'h1B3;
        15'h16CB: data = 12'h1B8;
        15'h16CC: data = 12'h1BD;
        15'h16CD: data = 12'h1C4;
        15'h16CE: data = 12'h1CA;
        15'h16CF: data = 12'h1CF;
        15'h16D0: data = 12'h1D0;
        15'h16D1: data = 12'h1DA;
        15'h16D2: data = 12'h1E2;
        15'h16D3: data = 12'h1EB;
        15'h16D4: data = 12'h1F9;
        15'h16D5: data = 12'h204;
        15'h16D6: data = 12'h211;
        15'h16D7: data = 12'h21C;
        15'h16D8: data = 12'h22D;
        15'h16D9: data = 12'h237;
        15'h16DA: data = 12'h247;
        15'h16DB: data = 12'h24F;
        15'h16DC: data = 12'h25E;
        15'h16DD: data = 12'h264;
        15'h16DE: data = 12'h271;
        15'h16DF: data = 12'h275;
        15'h16E0: data = 12'h285;
        15'h16E1: data = 12'h287;
        15'h16E2: data = 12'h295;
        15'h16E3: data = 12'h2A1;
        15'h16E4: data = 12'h2B0;
        15'h16E5: data = 12'h2BF;
        15'h16E6: data = 12'h2CD;
        15'h16E7: data = 12'h2DC;
        15'h16E8: data = 12'h2EC;
        15'h16E9: data = 12'h2FF;
        15'h16EA: data = 12'h310;
        15'h16EB: data = 12'h321;
        15'h16EC: data = 12'h332;
        15'h16ED: data = 12'h343;
        15'h16EE: data = 12'h356;
        15'h16EF: data = 12'h367;
        15'h16F0: data = 12'h377;
        15'h16F1: data = 12'h380;
        15'h16F2: data = 12'h397;
        15'h16F3: data = 12'h39D;
        15'h16F4: data = 12'h3B0;
        15'h16F5: data = 12'h3BC;
        15'h16F6: data = 12'h3C8;
        15'h16F7: data = 12'h3DC;
        15'h16F8: data = 12'h3EF;
        15'h16F9: data = 12'h400;
        15'h16FA: data = 12'h414;
        15'h16FB: data = 12'h425;
        15'h16FC: data = 12'h439;
        15'h16FD: data = 12'h450;
        15'h16FE: data = 12'h468;
        15'h16FF: data = 12'h47C;
        15'h1700: data = 12'h490;
        15'h1701: data = 12'h4A7;
        15'h1702: data = 12'h4B8;
        15'h1703: data = 12'h4D1;
        15'h1704: data = 12'h4E2;
        15'h1705: data = 12'h4F7;
        15'h1706: data = 12'h50D;
        15'h1707: data = 12'h51B;
        15'h1708: data = 12'h52F;
        15'h1709: data = 12'h542;
        15'h170A: data = 12'h558;
        15'h170B: data = 12'h569;
        15'h170C: data = 12'h578;
        15'h170D: data = 12'h58C;
        15'h170E: data = 12'h59E;
        15'h170F: data = 12'h5B2;
        15'h1710: data = 12'h5C7;
        15'h1711: data = 12'h5E0;
        15'h1712: data = 12'h5F7;
        15'h1713: data = 12'h612;
        15'h1714: data = 12'h628;
        15'h1715: data = 12'h63E;
        15'h1716: data = 12'h65A;
        15'h1717: data = 12'h675;
        15'h1718: data = 12'h68E;
        15'h1719: data = 12'h6A1;
        15'h171A: data = 12'h6B9;
        15'h171B: data = 12'h6D0;
        15'h171C: data = 12'h6E4;
        15'h171D: data = 12'h6F9;
        15'h171E: data = 12'h713;
        15'h171F: data = 12'h726;
        15'h1720: data = 12'h73D;
        15'h1721: data = 12'h74A;
        15'h1722: data = 12'h760;
        15'h1723: data = 12'h775;
        15'h1724: data = 12'h78E;
        15'h1725: data = 12'h7A0;
        15'h1726: data = 12'h7BB;
        15'h1727: data = 12'h7CF;
        15'h1728: data = 12'h7E3;
        15'h1729: data = 12'h7FD;
        15'h172A: data = 12'h06C;
        15'h172B: data = 12'h083;
        15'h172C: data = 12'h09D;
        15'h172D: data = 12'h0B0;
        15'h172E: data = 12'h0CB;
        15'h172F: data = 12'h0E6;
        15'h1730: data = 12'h100;
        15'h1731: data = 12'h110;
        15'h1732: data = 12'h12E;
        15'h1733: data = 12'h143;
        15'h1734: data = 12'h159;
        15'h1735: data = 12'h16D;
        15'h1736: data = 12'h182;
        15'h1737: data = 12'h19C;
        15'h1738: data = 12'h1B5;
        15'h1739: data = 12'h1C6;
        15'h173A: data = 12'h1DD;
        15'h173B: data = 12'h1F7;
        15'h173C: data = 12'h209;
        15'h173D: data = 12'h216;
        15'h173E: data = 12'h234;
        15'h173F: data = 12'h24B;
        15'h1740: data = 12'h263;
        15'h1741: data = 12'h272;
        15'h1742: data = 12'h289;
        15'h1743: data = 12'h2A5;
        15'h1744: data = 12'h2BC;
        15'h1745: data = 12'h2CE;
        15'h1746: data = 12'h2E8;
        15'h1747: data = 12'h2FE;
        15'h1748: data = 12'h31E;
        15'h1749: data = 12'h331;
        15'h174A: data = 12'h346;
        15'h174B: data = 12'h361;
        15'h174C: data = 12'h37A;
        15'h174D: data = 12'h394;
        15'h174E: data = 12'h3A8;
        15'h174F: data = 12'h3C3;
        15'h1750: data = 12'h3D9;
        15'h1751: data = 12'h3EF;
        15'h1752: data = 12'h3FF;
        15'h1753: data = 12'h414;
        15'h1754: data = 12'h42C;
        15'h1755: data = 12'h445;
        15'h1756: data = 12'h454;
        15'h1757: data = 12'h469;
        15'h1758: data = 12'h480;
        15'h1759: data = 12'h499;
        15'h175A: data = 12'h4AD;
        15'h175B: data = 12'h4C0;
        15'h175C: data = 12'h4CB;
        15'h175D: data = 12'h4DF;
        15'h175E: data = 12'h4F5;
        15'h175F: data = 12'h50A;
        15'h1760: data = 12'h515;
        15'h1761: data = 12'h528;
        15'h1762: data = 12'h53D;
        15'h1763: data = 12'h549;
        15'h1764: data = 12'h560;
        15'h1765: data = 12'h56E;
        15'h1766: data = 12'h583;
        15'h1767: data = 12'h595;
        15'h1768: data = 12'h5A6;
        15'h1769: data = 12'h5BA;
        15'h176A: data = 12'h5C3;
        15'h176B: data = 12'h5D5;
        15'h176C: data = 12'h5E8;
        15'h176D: data = 12'h5F9;
        15'h176E: data = 12'h60A;
        15'h176F: data = 12'h61B;
        15'h1770: data = 12'h62A;
        15'h1771: data = 12'h636;
        15'h1772: data = 12'h64B;
        15'h1773: data = 12'h660;
        15'h1774: data = 12'h66D;
        15'h1775: data = 12'h678;
        15'h1776: data = 12'h68C;
        15'h1777: data = 12'h69B;
        15'h1778: data = 12'h6AD;
        15'h1779: data = 12'h6BB;
        15'h177A: data = 12'h6CB;
        15'h177B: data = 12'h6D5;
        15'h177C: data = 12'h6E8;
        15'h177D: data = 12'h6F8;
        15'h177E: data = 12'h702;
        15'h177F: data = 12'h713;
        15'h1780: data = 12'h721;
        15'h1781: data = 12'h72F;
        15'h1782: data = 12'h737;
        15'h1783: data = 12'h741;
        15'h1784: data = 12'h74B;
        15'h1785: data = 12'h761;
        15'h1786: data = 12'h768;
        15'h1787: data = 12'h776;
        15'h1788: data = 12'h77E;
        15'h1789: data = 12'h78D;
        15'h178A: data = 12'h796;
        15'h178B: data = 12'h79C;
        15'h178C: data = 12'h7A3;
        15'h178D: data = 12'h7B1;
        15'h178E: data = 12'h7B9;
        15'h178F: data = 12'h7C2;
        15'h1790: data = 12'h7C6;
        15'h1791: data = 12'h7D2;
        15'h1792: data = 12'h7D9;
        15'h1793: data = 12'h7DE;
        15'h1794: data = 12'h7E6;
        15'h1795: data = 12'h7ED;
        15'h1796: data = 12'h7F3;
        15'h1797: data = 12'h7FA;
        15'h1798: data = 12'h804;
        15'h1799: data = 12'h801;
        15'h179A: data = 12'h808;
        15'h179B: data = 12'h80E;
        15'h179C: data = 12'h091;
        15'h179D: data = 12'h092;
        15'h179E: data = 12'h099;
        15'h179F: data = 12'h09C;
        15'h17A0: data = 12'h09F;
        15'h17A1: data = 12'h0A5;
        15'h17A2: data = 12'h0A4;
        15'h17A3: data = 12'h0AE;
        15'h17A4: data = 12'h0AA;
        15'h17A5: data = 12'h0AB;
        15'h17A6: data = 12'h0B4;
        15'h17A7: data = 12'h0B8;
        15'h17A8: data = 12'h0B9;
        15'h17A9: data = 12'h0B7;
        15'h17AA: data = 12'h0C0;
        15'h17AB: data = 12'h0C2;
        15'h17AC: data = 12'h0C7;
        15'h17AD: data = 12'h0CB;
        15'h17AE: data = 12'h0D1;
        15'h17AF: data = 12'h0D0;
        15'h17B0: data = 12'h0D4;
        15'h17B1: data = 12'h0CC;
        15'h17B2: data = 12'h0CD;
        15'h17B3: data = 12'h0CE;
        15'h17B4: data = 12'h0CD;
        15'h17B5: data = 12'h0CA;
        15'h17B6: data = 12'h0C1;
        15'h17B7: data = 12'h0BC;
        15'h17B8: data = 12'h0B0;
        15'h17B9: data = 12'h0AD;
        15'h17BA: data = 12'h0A6;
        15'h17BB: data = 12'h0A7;
        15'h17BC: data = 12'h0A8;
        15'h17BD: data = 12'h0AE;
        15'h17BE: data = 12'h0AA;
        15'h17BF: data = 12'h0A9;
        15'h17C0: data = 12'h0A7;
        15'h17C1: data = 12'h09F;
        15'h17C2: data = 12'h093;
        15'h17C3: data = 12'h089;
        15'h17C4: data = 12'h07A;
        15'h17C5: data = 12'h079;
        15'h17C6: data = 12'h06B;
        15'h17C7: data = 12'h06A;
        15'h17C8: data = 12'h066;
        15'h17C9: data = 12'h063;
        15'h17CA: data = 12'h061;
        15'h17CB: data = 12'h05B;
        15'h17CC: data = 12'h051;
        15'h17CD: data = 12'h000;
        15'h17CE: data = 12'h7B8;
        15'h17CF: data = 12'h7A8;
        15'h17D0: data = 12'h79F;
        15'h17D1: data = 12'h792;
        15'h17D2: data = 12'h78D;
        15'h17D3: data = 12'h78C;
        15'h17D4: data = 12'h77D;
        15'h17D5: data = 12'h772;
        15'h17D6: data = 12'h75F;
        15'h17D7: data = 12'h74E;
        15'h17D8: data = 12'h73B;
        15'h17D9: data = 12'h72E;
        15'h17DA: data = 12'h722;
        15'h17DB: data = 12'h717;
        15'h17DC: data = 12'h710;
        15'h17DD: data = 12'h70B;
        15'h17DE: data = 12'h6FD;
        15'h17DF: data = 12'h6EA;
        15'h17E0: data = 12'h6E0;
        15'h17E1: data = 12'h6CD;
        15'h17E2: data = 12'h6B8;
        15'h17E3: data = 12'h6A7;
        15'h17E4: data = 12'h693;
        15'h17E5: data = 12'h685;
        15'h17E6: data = 12'h676;
        15'h17E7: data = 12'h66A;
        15'h17E8: data = 12'h661;
        15'h17E9: data = 12'h655;
        15'h17EA: data = 12'h64A;
        15'h17EB: data = 12'h638;
        15'h17EC: data = 12'h62D;
        15'h17ED: data = 12'h615;
        15'h17EE: data = 12'h605;
        15'h17EF: data = 12'h5EF;
        15'h17F0: data = 12'h5D6;
        15'h17F1: data = 12'h5BF;
        15'h17F2: data = 12'h5B3;
        15'h17F3: data = 12'h5A3;
        15'h17F4: data = 12'h58C;
        15'h17F5: data = 12'h57E;
        15'h17F6: data = 12'h56A;
        15'h17F7: data = 12'h55A;
        15'h17F8: data = 12'h550;
        15'h17F9: data = 12'h540;
        15'h17FA: data = 12'h527;
        15'h17FB: data = 12'h51C;
        15'h17FC: data = 12'h506;
        15'h17FD: data = 12'h4F5;
        15'h17FE: data = 12'h4DB;
        15'h17FF: data = 12'h4CB;
        15'h1800: data = 12'h4B9;
        15'h1801: data = 12'h4A0;
        15'h1802: data = 12'h48B;
        15'h1803: data = 12'h472;
        15'h1804: data = 12'h459;
        15'h1805: data = 12'h444;
        15'h1806: data = 12'h430;
        15'h1807: data = 12'h415;
        15'h1808: data = 12'h400;
        15'h1809: data = 12'h3E8;
        15'h180A: data = 12'h3D6;
        15'h180B: data = 12'h3C0;
        15'h180C: data = 12'h3AA;
        15'h180D: data = 12'h38E;
        15'h180E: data = 12'h37C;
        15'h180F: data = 12'h366;
        15'h1810: data = 12'h351;
        15'h1811: data = 12'h33A;
        15'h1812: data = 12'h328;
        15'h1813: data = 12'h311;
        15'h1814: data = 12'h2F9;
        15'h1815: data = 12'h2E4;
        15'h1816: data = 12'h2D2;
        15'h1817: data = 12'h2BD;
        15'h1818: data = 12'h2A4;
        15'h1819: data = 12'h289;
        15'h181A: data = 12'h27A;
        15'h181B: data = 12'h262;
        15'h181C: data = 12'h247;
        15'h181D: data = 12'h232;
        15'h181E: data = 12'h217;
        15'h181F: data = 12'h205;
        15'h1820: data = 12'h1F2;
        15'h1821: data = 12'h1D8;
        15'h1822: data = 12'h1BF;
        15'h1823: data = 12'h1AA;
        15'h1824: data = 12'h191;
        15'h1825: data = 12'h17B;
        15'h1826: data = 12'h163;
        15'h1827: data = 12'h14E;
        15'h1828: data = 12'h131;
        15'h1829: data = 12'h11B;
        15'h182A: data = 12'h109;
        15'h182B: data = 12'h0F0;
        15'h182C: data = 12'h0DA;
        15'h182D: data = 12'h0BF;
        15'h182E: data = 12'h0A5;
        15'h182F: data = 12'h090;
        15'h1830: data = 12'h080;
        15'h1831: data = 12'h063;
        15'h1832: data = 12'h04F;
        15'h1833: data = 12'h7E3;
        15'h1834: data = 12'h7CE;
        15'h1835: data = 12'h7B8;
        15'h1836: data = 12'h7A4;
        15'h1837: data = 12'h78B;
        15'h1838: data = 12'h776;
        15'h1839: data = 12'h75E;
        15'h183A: data = 12'h74C;
        15'h183B: data = 12'h735;
        15'h183C: data = 12'h71D;
        15'h183D: data = 12'h706;
        15'h183E: data = 12'h6EE;
        15'h183F: data = 12'h6DB;
        15'h1840: data = 12'h6C5;
        15'h1841: data = 12'h6AC;
        15'h1842: data = 12'h698;
        15'h1843: data = 12'h685;
        15'h1844: data = 12'h668;
        15'h1845: data = 12'h657;
        15'h1846: data = 12'h63C;
        15'h1847: data = 12'h62F;
        15'h1848: data = 12'h618;
        15'h1849: data = 12'h600;
        15'h184A: data = 12'h5E7;
        15'h184B: data = 12'h5D1;
        15'h184C: data = 12'h5C5;
        15'h184D: data = 12'h5A2;
        15'h184E: data = 12'h58F;
        15'h184F: data = 12'h578;
        15'h1850: data = 12'h565;
        15'h1851: data = 12'h552;
        15'h1852: data = 12'h53B;
        15'h1853: data = 12'h522;
        15'h1854: data = 12'h511;
        15'h1855: data = 12'h4F7;
        15'h1856: data = 12'h4E0;
        15'h1857: data = 12'h4CD;
        15'h1858: data = 12'h4B7;
        15'h1859: data = 12'h4A5;
        15'h185A: data = 12'h492;
        15'h185B: data = 12'h47C;
        15'h185C: data = 12'h466;
        15'h185D: data = 12'h452;
        15'h185E: data = 12'h443;
        15'h185F: data = 12'h436;
        15'h1860: data = 12'h420;
        15'h1861: data = 12'h414;
        15'h1862: data = 12'h402;
        15'h1863: data = 12'h3F5;
        15'h1864: data = 12'h3E8;
        15'h1865: data = 12'h3D0;
        15'h1866: data = 12'h3C0;
        15'h1867: data = 12'h3B5;
        15'h1868: data = 12'h39E;
        15'h1869: data = 12'h393;
        15'h186A: data = 12'h37E;
        15'h186B: data = 12'h36D;
        15'h186C: data = 12'h35D;
        15'h186D: data = 12'h349;
        15'h186E: data = 12'h336;
        15'h186F: data = 12'h320;
        15'h1870: data = 12'h30E;
        15'h1871: data = 12'h2FF;
        15'h1872: data = 12'h2F0;
        15'h1873: data = 12'h2DD;
        15'h1874: data = 12'h2D2;
        15'h1875: data = 12'h2C9;
        15'h1876: data = 12'h2BF;
        15'h1877: data = 12'h2B0;
        15'h1878: data = 12'h2A9;
        15'h1879: data = 12'h29F;
        15'h187A: data = 12'h295;
        15'h187B: data = 12'h288;
        15'h187C: data = 12'h281;
        15'h187D: data = 12'h26D;
        15'h187E: data = 12'h265;
        15'h187F: data = 12'h250;
        15'h1880: data = 12'h247;
        15'h1881: data = 12'h233;
        15'h1882: data = 12'h226;
        15'h1883: data = 12'h218;
        15'h1884: data = 12'h210;
        15'h1885: data = 12'h208;
        15'h1886: data = 12'h202;
        15'h1887: data = 12'h1F3;
        15'h1888: data = 12'h1ED;
        15'h1889: data = 12'h1E8;
        15'h188A: data = 12'h1E6;
        15'h188B: data = 12'h1E6;
        15'h188C: data = 12'h1D8;
        15'h188D: data = 12'h1CE;
        15'h188E: data = 12'h1C6;
        15'h188F: data = 12'h1C3;
        15'h1890: data = 12'h1B7;
        15'h1891: data = 12'h1AB;
        15'h1892: data = 12'h19F;
        15'h1893: data = 12'h195;
        15'h1894: data = 12'h193;
        15'h1895: data = 12'h189;
        15'h1896: data = 12'h185;
        15'h1897: data = 12'h185;
        15'h1898: data = 12'h182;
        15'h1899: data = 12'h181;
        15'h189A: data = 12'h182;
        15'h189B: data = 12'h17F;
        15'h189C: data = 12'h17C;
        15'h189D: data = 12'h174;
        15'h189E: data = 12'h177;
        15'h189F: data = 12'h173;
        15'h18A0: data = 12'h169;
        15'h18A1: data = 12'h163;
        15'h18A2: data = 12'h163;
        15'h18A3: data = 12'h160;
        15'h18A4: data = 12'h157;
        15'h18A5: data = 12'h154;
        15'h18A6: data = 12'h157;
        15'h18A7: data = 12'h159;
        15'h18A8: data = 12'h15D;
        15'h18A9: data = 12'h164;
        15'h18AA: data = 12'h164;
        15'h18AB: data = 12'h16C;
        15'h18AC: data = 12'h170;
        15'h18AD: data = 12'h16D;
        15'h18AE: data = 12'h16C;
        15'h18AF: data = 12'h16D;
        15'h18B0: data = 12'h170;
        15'h18B1: data = 12'h16F;
        15'h18B2: data = 12'h16D;
        15'h18B3: data = 12'h16F;
        15'h18B4: data = 12'h16D;
        15'h18B5: data = 12'h177;
        15'h18B6: data = 12'h17E;
        15'h18B7: data = 12'h181;
        15'h18B8: data = 12'h189;
        15'h18B9: data = 12'h18B;
        15'h18BA: data = 12'h19C;
        15'h18BB: data = 12'h1A1;
        15'h18BC: data = 12'h1AD;
        15'h18BD: data = 12'h1B3;
        15'h18BE: data = 12'h1B1;
        15'h18BF: data = 12'h1BA;
        15'h18C0: data = 12'h1C2;
        15'h18C1: data = 12'h1C4;
        15'h18C2: data = 12'h1C8;
        15'h18C3: data = 12'h1D0;
        15'h18C4: data = 12'h1D2;
        15'h18C5: data = 12'h1D9;
        15'h18C6: data = 12'h1DF;
        15'h18C7: data = 12'h1EF;
        15'h18C8: data = 12'h1FA;
        15'h18C9: data = 12'h206;
        15'h18CA: data = 12'h214;
        15'h18CB: data = 12'h219;
        15'h18CC: data = 12'h22D;
        15'h18CD: data = 12'h236;
        15'h18CE: data = 12'h247;
        15'h18CF: data = 12'h24F;
        15'h18D0: data = 12'h260;
        15'h18D1: data = 12'h266;
        15'h18D2: data = 12'h276;
        15'h18D3: data = 12'h277;
        15'h18D4: data = 12'h284;
        15'h18D5: data = 12'h28B;
        15'h18D6: data = 12'h293;
        15'h18D7: data = 12'h2A1;
        15'h18D8: data = 12'h2B0;
        15'h18D9: data = 12'h2BD;
        15'h18DA: data = 12'h2CD;
        15'h18DB: data = 12'h2D9;
        15'h18DC: data = 12'h2E9;
        15'h18DD: data = 12'h2FF;
        15'h18DE: data = 12'h313;
        15'h18DF: data = 12'h325;
        15'h18E0: data = 12'h337;
        15'h18E1: data = 12'h344;
        15'h18E2: data = 12'h357;
        15'h18E3: data = 12'h367;
        15'h18E4: data = 12'h375;
        15'h18E5: data = 12'h380;
        15'h18E6: data = 12'h396;
        15'h18E7: data = 12'h39F;
        15'h18E8: data = 12'h3AF;
        15'h18E9: data = 12'h3BB;
        15'h18EA: data = 12'h3C8;
        15'h18EB: data = 12'h3E0;
        15'h18EC: data = 12'h3EF;
        15'h18ED: data = 12'h3FC;
        15'h18EE: data = 12'h415;
        15'h18EF: data = 12'h428;
        15'h18F0: data = 12'h436;
        15'h18F1: data = 12'h452;
        15'h18F2: data = 12'h465;
        15'h18F3: data = 12'h47E;
        15'h18F4: data = 12'h490;
        15'h18F5: data = 12'h4AA;
        15'h18F6: data = 12'h4BA;
        15'h18F7: data = 12'h4D2;
        15'h18F8: data = 12'h4E1;
        15'h18F9: data = 12'h4F5;
        15'h18FA: data = 12'h50A;
        15'h18FB: data = 12'h51D;
        15'h18FC: data = 12'h52F;
        15'h18FD: data = 12'h543;
        15'h18FE: data = 12'h557;
        15'h18FF: data = 12'h565;
        15'h1900: data = 12'h578;
        15'h1901: data = 12'h58A;
        15'h1902: data = 12'h59E;
        15'h1903: data = 12'h5B0;
        15'h1904: data = 12'h5CA;
        15'h1905: data = 12'h5E2;
        15'h1906: data = 12'h5F8;
        15'h1907: data = 12'h615;
        15'h1908: data = 12'h62A;
        15'h1909: data = 12'h643;
        15'h190A: data = 12'h65C;
        15'h190B: data = 12'h672;
        15'h190C: data = 12'h68D;
        15'h190D: data = 12'h6A2;
        15'h190E: data = 12'h6B7;
        15'h190F: data = 12'h6CF;
        15'h1910: data = 12'h6E0;
        15'h1911: data = 12'h6FA;
        15'h1912: data = 12'h70F;
        15'h1913: data = 12'h722;
        15'h1914: data = 12'h73A;
        15'h1915: data = 12'h74B;
        15'h1916: data = 12'h75E;
        15'h1917: data = 12'h776;
        15'h1918: data = 12'h78D;
        15'h1919: data = 12'h7A2;
        15'h191A: data = 12'h7B7;
        15'h191B: data = 12'h7D2;
        15'h191C: data = 12'h7E8;
        15'h191D: data = 12'h7FF;
        15'h191E: data = 12'h12A;
        15'h191F: data = 12'h087;
        15'h1920: data = 12'h09E;
        15'h1921: data = 12'h0B2;
        15'h1922: data = 12'h0CE;
        15'h1923: data = 12'h0E8;
        15'h1924: data = 12'h102;
        15'h1925: data = 12'h113;
        15'h1926: data = 12'h12E;
        15'h1927: data = 12'h144;
        15'h1928: data = 12'h159;
        15'h1929: data = 12'h170;
        15'h192A: data = 12'h183;
        15'h192B: data = 12'h19D;
        15'h192C: data = 12'h1B5;
        15'h192D: data = 12'h1C1;
        15'h192E: data = 12'h1D8;
        15'h192F: data = 12'h1F3;
        15'h1930: data = 12'h208;
        15'h1931: data = 12'h215;
        15'h1932: data = 12'h231;
        15'h1933: data = 12'h24C;
        15'h1934: data = 12'h25E;
        15'h1935: data = 12'h275;
        15'h1936: data = 12'h287;
        15'h1937: data = 12'h2A3;
        15'h1938: data = 12'h2BE;
        15'h1939: data = 12'h2CF;
        15'h193A: data = 12'h2E9;
        15'h193B: data = 12'h300;
        15'h193C: data = 12'h31E;
        15'h193D: data = 12'h330;
        15'h193E: data = 12'h348;
        15'h193F: data = 12'h364;
        15'h1940: data = 12'h37A;
        15'h1941: data = 12'h398;
        15'h1942: data = 12'h3A8;
        15'h1943: data = 12'h3C5;
        15'h1944: data = 12'h3DB;
        15'h1945: data = 12'h3EE;
        15'h1946: data = 12'h3FE;
        15'h1947: data = 12'h415;
        15'h1948: data = 12'h430;
        15'h1949: data = 12'h447;
        15'h194A: data = 12'h452;
        15'h194B: data = 12'h46D;
        15'h194C: data = 12'h482;
        15'h194D: data = 12'h495;
        15'h194E: data = 12'h4AA;
        15'h194F: data = 12'h4BD;
        15'h1950: data = 12'h4C9;
        15'h1951: data = 12'h4E0;
        15'h1952: data = 12'h4F4;
        15'h1953: data = 12'h50A;
        15'h1954: data = 12'h514;
        15'h1955: data = 12'h529;
        15'h1956: data = 12'h53E;
        15'h1957: data = 12'h548;
        15'h1958: data = 12'h561;
        15'h1959: data = 12'h56E;
        15'h195A: data = 12'h583;
        15'h195B: data = 12'h594;
        15'h195C: data = 12'h5A4;
        15'h195D: data = 12'h5BB;
        15'h195E: data = 12'h5C2;
        15'h195F: data = 12'h5D3;
        15'h1960: data = 12'h5EB;
        15'h1961: data = 12'h5FA;
        15'h1962: data = 12'h60B;
        15'h1963: data = 12'h619;
        15'h1964: data = 12'h62A;
        15'h1965: data = 12'h637;
        15'h1966: data = 12'h64D;
        15'h1967: data = 12'h65F;
        15'h1968: data = 12'h671;
        15'h1969: data = 12'h67C;
        15'h196A: data = 12'h690;
        15'h196B: data = 12'h6A2;
        15'h196C: data = 12'h6AC;
        15'h196D: data = 12'h6BB;
        15'h196E: data = 12'h6CC;
        15'h196F: data = 12'h6D8;
        15'h1970: data = 12'h6EA;
        15'h1971: data = 12'h6FA;
        15'h1972: data = 12'h706;
        15'h1973: data = 12'h712;
        15'h1974: data = 12'h725;
        15'h1975: data = 12'h735;
        15'h1976: data = 12'h736;
        15'h1977: data = 12'h741;
        15'h1978: data = 12'h752;
        15'h1979: data = 12'h75F;
        15'h197A: data = 12'h76A;
        15'h197B: data = 12'h776;
        15'h197C: data = 12'h77D;
        15'h197D: data = 12'h790;
        15'h197E: data = 12'h79A;
        15'h197F: data = 12'h79D;
        15'h1980: data = 12'h7A4;
        15'h1981: data = 12'h7B0;
        15'h1982: data = 12'h7BB;
        15'h1983: data = 12'h7C2;
        15'h1984: data = 12'h7C9;
        15'h1985: data = 12'h7CE;
        15'h1986: data = 12'h7D6;
        15'h1987: data = 12'h7E0;
        15'h1988: data = 12'h7E9;
        15'h1989: data = 12'h7EC;
        15'h198A: data = 12'h7F4;
        15'h198B: data = 12'h7FA;
        15'h198C: data = 12'h802;
        15'h198D: data = 12'h804;
        15'h198E: data = 12'h80A;
        15'h198F: data = 12'h079;
        15'h1990: data = 12'h091;
        15'h1991: data = 12'h092;
        15'h1992: data = 12'h099;
        15'h1993: data = 12'h09E;
        15'h1994: data = 12'h09E;
        15'h1995: data = 12'h0A7;
        15'h1996: data = 12'h0A8;
        15'h1997: data = 12'h0AE;
        15'h1998: data = 12'h0B1;
        15'h1999: data = 12'h0AF;
        15'h199A: data = 12'h0B9;
        15'h199B: data = 12'h0B9;
        15'h199C: data = 12'h0BA;
        15'h199D: data = 12'h0BD;
        15'h199E: data = 12'h0C1;
        15'h199F: data = 12'h0C8;
        15'h19A0: data = 12'h0CA;
        15'h19A1: data = 12'h0CD;
        15'h19A2: data = 12'h0D5;
        15'h19A3: data = 12'h0D5;
        15'h19A4: data = 12'h0D5;
        15'h19A5: data = 12'h0CB;
        15'h19A6: data = 12'h0CE;
        15'h19A7: data = 12'h0CC;
        15'h19A8: data = 12'h0CA;
        15'h19A9: data = 12'h0C8;
        15'h19AA: data = 12'h0BC;
        15'h19AB: data = 12'h0B5;
        15'h19AC: data = 12'h0AC;
        15'h19AD: data = 12'h0AC;
        15'h19AE: data = 12'h0A8;
        15'h19AF: data = 12'h0A9;
        15'h19B0: data = 12'h0AB;
        15'h19B1: data = 12'h0AD;
        15'h19B2: data = 12'h0AA;
        15'h19B3: data = 12'h0A7;
        15'h19B4: data = 12'h0A6;
        15'h19B5: data = 12'h09B;
        15'h19B6: data = 12'h092;
        15'h19B7: data = 12'h07D;
        15'h19B8: data = 12'h073;
        15'h19B9: data = 12'h073;
        15'h19BA: data = 12'h06D;
        15'h19BB: data = 12'h06C;
        15'h19BC: data = 12'h06B;
        15'h19BD: data = 12'h068;
        15'h19BE: data = 12'h060;
        15'h19BF: data = 12'h058;
        15'h19C0: data = 12'h047;
        15'h19C1: data = 12'h7BE;
        15'h19C2: data = 12'h7B2;
        15'h19C3: data = 12'h7A6;
        15'h19C4: data = 12'h7A2;
        15'h19C5: data = 12'h79D;
        15'h19C6: data = 12'h793;
        15'h19C7: data = 12'h78D;
        15'h19C8: data = 12'h779;
        15'h19C9: data = 12'h770;
        15'h19CA: data = 12'h756;
        15'h19CB: data = 12'h746;
        15'h19CC: data = 12'h735;
        15'h19CD: data = 12'h72B;
        15'h19CE: data = 12'h724;
        15'h19CF: data = 12'h71D;
        15'h19D0: data = 12'h715;
        15'h19D1: data = 12'h70B;
        15'h19D2: data = 12'h6F8;
        15'h19D3: data = 12'h6E9;
        15'h19D4: data = 12'h6DB;
        15'h19D5: data = 12'h6C7;
        15'h19D6: data = 12'h6B1;
        15'h19D7: data = 12'h6A0;
        15'h19D8: data = 12'h698;
        15'h19D9: data = 12'h687;
        15'h19DA: data = 12'h67D;
        15'h19DB: data = 12'h672;
        15'h19DC: data = 12'h665;
        15'h19DD: data = 12'h656;
        15'h19DE: data = 12'h647;
        15'h19DF: data = 12'h635;
        15'h19E0: data = 12'h629;
        15'h19E1: data = 12'h60E;
        15'h19E2: data = 12'h5FC;
        15'h19E3: data = 12'h5E9;
        15'h19E4: data = 12'h5CF;
        15'h19E5: data = 12'h5BC;
        15'h19E6: data = 12'h5B1;
        15'h19E7: data = 12'h5A4;
        15'h19E8: data = 12'h590;
        15'h19E9: data = 12'h581;
        15'h19EA: data = 12'h56F;
        15'h19EB: data = 12'h567;
        15'h19EC: data = 12'h554;
        15'h19ED: data = 12'h544;
        15'h19EE: data = 12'h52C;
        15'h19EF: data = 12'h51C;
        15'h19F0: data = 12'h506;
        15'h19F1: data = 12'h4F2;
        15'h19F2: data = 12'h4DB;
        15'h19F3: data = 12'h4C2;
        15'h19F4: data = 12'h4AF;
        15'h19F5: data = 12'h497;
        15'h19F6: data = 12'h481;
        15'h19F7: data = 12'h469;
        15'h19F8: data = 12'h455;
        15'h19F9: data = 12'h442;
        15'h19FA: data = 12'h42C;
        15'h19FB: data = 12'h414;
        15'h19FC: data = 12'h3FD;
        15'h19FD: data = 12'h3E8;
        15'h19FE: data = 12'h3D4;
        15'h19FF: data = 12'h3C3;
        15'h1A00: data = 12'h3AE;
        15'h1A01: data = 12'h392;
        15'h1A02: data = 12'h384;
        15'h1A03: data = 12'h36C;
        15'h1A04: data = 12'h357;
        15'h1A05: data = 12'h33D;
        15'h1A06: data = 12'h32D;
        15'h1A07: data = 12'h31B;
        15'h1A08: data = 12'h300;
        15'h1A09: data = 12'h2EB;
        15'h1A0A: data = 12'h2D8;
        15'h1A0B: data = 12'h2C2;
        15'h1A0C: data = 12'h2AD;
        15'h1A0D: data = 12'h28F;
        15'h1A0E: data = 12'h280;
        15'h1A0F: data = 12'h268;
        15'h1A10: data = 12'h24B;
        15'h1A11: data = 12'h237;
        15'h1A12: data = 12'h21E;
        15'h1A13: data = 12'h206;
        15'h1A14: data = 12'h1F6;
        15'h1A15: data = 12'h1DA;
        15'h1A16: data = 12'h1C1;
        15'h1A17: data = 12'h1A9;
        15'h1A18: data = 12'h194;
        15'h1A19: data = 12'h181;
        15'h1A1A: data = 12'h168;
        15'h1A1B: data = 12'h14D;
        15'h1A1C: data = 12'h13A;
        15'h1A1D: data = 12'h11E;
        15'h1A1E: data = 12'h10B;
        15'h1A1F: data = 12'h0F5;
        15'h1A20: data = 12'h0DB;
        15'h1A21: data = 12'h0C2;
        15'h1A22: data = 12'h0A9;
        15'h1A23: data = 12'h093;
        15'h1A24: data = 12'h082;
        15'h1A25: data = 12'h067;
        15'h1A26: data = 12'h04C;
        15'h1A27: data = 12'h7E0;
        15'h1A28: data = 12'h7D0;
        15'h1A29: data = 12'h7BC;
        15'h1A2A: data = 12'h7A5;
        15'h1A2B: data = 12'h78D;
        15'h1A2C: data = 12'h775;
        15'h1A2D: data = 12'h760;
        15'h1A2E: data = 12'h74B;
        15'h1A2F: data = 12'h736;
        15'h1A30: data = 12'h71E;
        15'h1A31: data = 12'h705;
        15'h1A32: data = 12'h6F0;
        15'h1A33: data = 12'h6D8;
        15'h1A34: data = 12'h6C4;
        15'h1A35: data = 12'h6AE;
        15'h1A36: data = 12'h698;
        15'h1A37: data = 12'h682;
        15'h1A38: data = 12'h669;
        15'h1A39: data = 12'h658;
        15'h1A3A: data = 12'h639;
        15'h1A3B: data = 12'h62C;
        15'h1A3C: data = 12'h616;
        15'h1A3D: data = 12'h5FB;
        15'h1A3E: data = 12'h5E7;
        15'h1A3F: data = 12'h5CF;
        15'h1A40: data = 12'h5C0;
        15'h1A41: data = 12'h5A2;
        15'h1A42: data = 12'h58B;
        15'h1A43: data = 12'h578;
        15'h1A44: data = 12'h562;
        15'h1A45: data = 12'h54C;
        15'h1A46: data = 12'h534;
        15'h1A47: data = 12'h51B;
        15'h1A48: data = 12'h50F;
        15'h1A49: data = 12'h4F5;
        15'h1A4A: data = 12'h4DC;
        15'h1A4B: data = 12'h4CB;
        15'h1A4C: data = 12'h4B8;
        15'h1A4D: data = 12'h4A5;
        15'h1A4E: data = 12'h491;
        15'h1A4F: data = 12'h47E;
        15'h1A50: data = 12'h46C;
        15'h1A51: data = 12'h457;
        15'h1A52: data = 12'h449;
        15'h1A53: data = 12'h43C;
        15'h1A54: data = 12'h428;
        15'h1A55: data = 12'h419;
        15'h1A56: data = 12'h404;
        15'h1A57: data = 12'h3FA;
        15'h1A58: data = 12'h3E8;
        15'h1A59: data = 12'h3D4;
        15'h1A5A: data = 12'h3C1;
        15'h1A5B: data = 12'h3B2;
        15'h1A5C: data = 12'h39E;
        15'h1A5D: data = 12'h392;
        15'h1A5E: data = 12'h379;
        15'h1A5F: data = 12'h366;
        15'h1A60: data = 12'h352;
        15'h1A61: data = 12'h343;
        15'h1A62: data = 12'h333;
        15'h1A63: data = 12'h31F;
        15'h1A64: data = 12'h30F;
        15'h1A65: data = 12'h2FF;
        15'h1A66: data = 12'h2F2;
        15'h1A67: data = 12'h2E4;
        15'h1A68: data = 12'h2D4;
        15'h1A69: data = 12'h2CF;
        15'h1A6A: data = 12'h2C5;
        15'h1A6B: data = 12'h2B7;
        15'h1A6C: data = 12'h2AC;
        15'h1A6D: data = 12'h2A2;
        15'h1A6E: data = 12'h295;
        15'h1A6F: data = 12'h284;
        15'h1A70: data = 12'h27F;
        15'h1A71: data = 12'h26E;
        15'h1A72: data = 12'h25E;
        15'h1A73: data = 12'h253;
        15'h1A74: data = 12'h243;
        15'h1A75: data = 12'h22D;
        15'h1A76: data = 12'h227;
        15'h1A77: data = 12'h215;
        15'h1A78: data = 12'h20D;
        15'h1A79: data = 12'h20A;
        15'h1A7A: data = 12'h202;
        15'h1A7B: data = 12'h1F7;
        15'h1A7C: data = 12'h1F3;
        15'h1A7D: data = 12'h1ED;
        15'h1A7E: data = 12'h1EB;
        15'h1A7F: data = 12'h1E3;
        15'h1A80: data = 12'h1D7;
        15'h1A81: data = 12'h1CB;
        15'h1A82: data = 12'h1C7;
        15'h1A83: data = 12'h1BE;
        15'h1A84: data = 12'h1B5;
        15'h1A85: data = 12'h1A6;
        15'h1A86: data = 12'h19D;
        15'h1A87: data = 12'h198;
        15'h1A88: data = 12'h194;
        15'h1A89: data = 12'h18D;
        15'h1A8A: data = 12'h185;
        15'h1A8B: data = 12'h187;
        15'h1A8C: data = 12'h188;
        15'h1A8D: data = 12'h187;
        15'h1A8E: data = 12'h184;
        15'h1A8F: data = 12'h181;
        15'h1A90: data = 12'h17D;
        15'h1A91: data = 12'h179;
        15'h1A92: data = 12'h175;
        15'h1A93: data = 12'h171;
        15'h1A94: data = 12'h165;
        15'h1A95: data = 12'h162;
        15'h1A96: data = 12'h15F;
        15'h1A97: data = 12'h15E;
        15'h1A98: data = 12'h155;
        15'h1A99: data = 12'h158;
        15'h1A9A: data = 12'h157;
        15'h1A9B: data = 12'h15C;
        15'h1A9C: data = 12'h160;
        15'h1A9D: data = 12'h163;
        15'h1A9E: data = 12'h169;
        15'h1A9F: data = 12'h171;
        15'h1AA0: data = 12'h171;
        15'h1AA1: data = 12'h16D;
        15'h1AA2: data = 12'h16A;
        15'h1AA3: data = 12'h16B;
        15'h1AA4: data = 12'h16D;
        15'h1AA5: data = 12'h16A;
        15'h1AA6: data = 12'h168;
        15'h1AA7: data = 12'h16E;
        15'h1AA8: data = 12'h16C;
        15'h1AA9: data = 12'h174;
        15'h1AAA: data = 12'h17D;
        15'h1AAB: data = 12'h17F;
        15'h1AAC: data = 12'h18D;
        15'h1AAD: data = 12'h190;
        15'h1AAE: data = 12'h19C;
        15'h1AAF: data = 12'h1A7;
        15'h1AB0: data = 12'h1B0;
        15'h1AB1: data = 12'h1B6;
        15'h1AB2: data = 12'h1B8;
        15'h1AB3: data = 12'h1BA;
        15'h1AB4: data = 12'h1BE;
        15'h1AB5: data = 12'h1C1;
        15'h1AB6: data = 12'h1C8;
        15'h1AB7: data = 12'h1C7;
        15'h1AB8: data = 12'h1D1;
        15'h1AB9: data = 12'h1D7;
        15'h1ABA: data = 12'h1E3;
        15'h1ABB: data = 12'h1ED;
        15'h1ABC: data = 12'h1FC;
        15'h1ABD: data = 12'h20A;
        15'h1ABE: data = 12'h216;
        15'h1ABF: data = 12'h220;
        15'h1AC0: data = 12'h231;
        15'h1AC1: data = 12'h239;
        15'h1AC2: data = 12'h249;
        15'h1AC3: data = 12'h24F;
        15'h1AC4: data = 12'h25D;
        15'h1AC5: data = 12'h261;
        15'h1AC6: data = 12'h271;
        15'h1AC7: data = 12'h270;
        15'h1AC8: data = 12'h280;
        15'h1AC9: data = 12'h288;
        15'h1ACA: data = 12'h292;
        15'h1ACB: data = 12'h2A3;
        15'h1ACC: data = 12'h2B2;
        15'h1ACD: data = 12'h2C0;
        15'h1ACE: data = 12'h2D1;
        15'h1ACF: data = 12'h2DD;
        15'h1AD0: data = 12'h2EF;
        15'h1AD1: data = 12'h302;
        15'h1AD2: data = 12'h315;
        15'h1AD3: data = 12'h325;
        15'h1AD4: data = 12'h33A;
        15'h1AD5: data = 12'h346;
        15'h1AD6: data = 12'h357;
        15'h1AD7: data = 12'h367;
        15'h1AD8: data = 12'h372;
        15'h1AD9: data = 12'h37E;
        15'h1ADA: data = 12'h390;
        15'h1ADB: data = 12'h398;
        15'h1ADC: data = 12'h3AD;
        15'h1ADD: data = 12'h3B8;
        15'h1ADE: data = 12'h3C9;
        15'h1ADF: data = 12'h3DD;
        15'h1AE0: data = 12'h3ED;
        15'h1AE1: data = 12'h3FD;
        15'h1AE2: data = 12'h412;
        15'h1AE3: data = 12'h429;
        15'h1AE4: data = 12'h43E;
        15'h1AE5: data = 12'h454;
        15'h1AE6: data = 12'h469;
        15'h1AE7: data = 12'h480;
        15'h1AE8: data = 12'h492;
        15'h1AE9: data = 12'h4A8;
        15'h1AEA: data = 12'h4B6;
        15'h1AEB: data = 12'h4D1;
        15'h1AEC: data = 12'h4E3;
        15'h1AED: data = 12'h4F7;
        15'h1AEE: data = 12'h50A;
        15'h1AEF: data = 12'h51A;
        15'h1AF0: data = 12'h52E;
        15'h1AF1: data = 12'h542;
        15'h1AF2: data = 12'h557;
        15'h1AF3: data = 12'h565;
        15'h1AF4: data = 12'h573;
        15'h1AF5: data = 12'h58C;
        15'h1AF6: data = 12'h59D;
        15'h1AF7: data = 12'h5B7;
        15'h1AF8: data = 12'h5CD;
        15'h1AF9: data = 12'h5E3;
        15'h1AFA: data = 12'h600;
        15'h1AFB: data = 12'h616;
        15'h1AFC: data = 12'h62C;
        15'h1AFD: data = 12'h643;
        15'h1AFE: data = 12'h662;
        15'h1AFF: data = 12'h677;
        15'h1B00: data = 12'h693;
        15'h1B01: data = 12'h6A1;
        15'h1B02: data = 12'h6B9;
        15'h1B03: data = 12'h6CF;
        15'h1B04: data = 12'h6E3;
        15'h1B05: data = 12'h6FA;
        15'h1B06: data = 12'h711;
        15'h1B07: data = 12'h724;
        15'h1B08: data = 12'h734;
        15'h1B09: data = 12'h748;
        15'h1B0A: data = 12'h75E;
        15'h1B0B: data = 12'h776;
        15'h1B0C: data = 12'h78E;
        15'h1B0D: data = 12'h79E;
        15'h1B0E: data = 12'h7B6;
        15'h1B0F: data = 12'h7D0;
        15'h1B10: data = 12'h7E6;
        15'h1B11: data = 12'h800;
        15'h1B12: data = 12'h06E;
        15'h1B13: data = 12'h087;
        15'h1B14: data = 12'h09C;
        15'h1B15: data = 12'h0B2;
        15'h1B16: data = 12'h0D1;
        15'h1B17: data = 12'h0EA;
        15'h1B18: data = 12'h101;
        15'h1B19: data = 12'h116;
        15'h1B1A: data = 12'h12E;
        15'h1B1B: data = 12'h142;
        15'h1B1C: data = 12'h157;
        15'h1B1D: data = 12'h16E;
        15'h1B1E: data = 12'h183;
        15'h1B1F: data = 12'h19C;
        15'h1B20: data = 12'h1B4;
        15'h1B21: data = 12'h1C0;
        15'h1B22: data = 12'h1DC;
        15'h1B23: data = 12'h1EF;
        15'h1B24: data = 12'h208;
        15'h1B25: data = 12'h219;
        15'h1B26: data = 12'h230;
        15'h1B27: data = 12'h24B;
        15'h1B28: data = 12'h25F;
        15'h1B29: data = 12'h271;
        15'h1B2A: data = 12'h28C;
        15'h1B2B: data = 12'h2A5;
        15'h1B2C: data = 12'h2BC;
        15'h1B2D: data = 12'h2D1;
        15'h1B2E: data = 12'h2ED;
        15'h1B2F: data = 12'h303;
        15'h1B30: data = 12'h321;
        15'h1B31: data = 12'h333;
        15'h1B32: data = 12'h34B;
        15'h1B33: data = 12'h365;
        15'h1B34: data = 12'h37C;
        15'h1B35: data = 12'h395;
        15'h1B36: data = 12'h3AA;
        15'h1B37: data = 12'h3C3;
        15'h1B38: data = 12'h3DC;
        15'h1B39: data = 12'h3F0;
        15'h1B3A: data = 12'h403;
        15'h1B3B: data = 12'h41A;
        15'h1B3C: data = 12'h42D;
        15'h1B3D: data = 12'h446;
        15'h1B3E: data = 12'h456;
        15'h1B3F: data = 12'h46A;
        15'h1B40: data = 12'h483;
        15'h1B41: data = 12'h496;
        15'h1B42: data = 12'h4AC;
        15'h1B43: data = 12'h4BE;
        15'h1B44: data = 12'h4C9;
        15'h1B45: data = 12'h4E0;
        15'h1B46: data = 12'h4F7;
        15'h1B47: data = 12'h50B;
        15'h1B48: data = 12'h517;
        15'h1B49: data = 12'h528;
        15'h1B4A: data = 12'h53F;
        15'h1B4B: data = 12'h54A;
        15'h1B4C: data = 12'h561;
        15'h1B4D: data = 12'h56D;
        15'h1B4E: data = 12'h584;
        15'h1B4F: data = 12'h593;
        15'h1B50: data = 12'h5A5;
        15'h1B51: data = 12'h5BA;
        15'h1B52: data = 12'h5C2;
        15'h1B53: data = 12'h5D4;
        15'h1B54: data = 12'h5ED;
        15'h1B55: data = 12'h5FD;
        15'h1B56: data = 12'h60E;
        15'h1B57: data = 12'h619;
        15'h1B58: data = 12'h62A;
        15'h1B59: data = 12'h636;
        15'h1B5A: data = 12'h64E;
        15'h1B5B: data = 12'h65D;
        15'h1B5C: data = 12'h670;
        15'h1B5D: data = 12'h67D;
        15'h1B5E: data = 12'h691;
        15'h1B5F: data = 12'h6A1;
        15'h1B60: data = 12'h6AF;
        15'h1B61: data = 12'h6C1;
        15'h1B62: data = 12'h6CD;
        15'h1B63: data = 12'h6D8;
        15'h1B64: data = 12'h6E8;
        15'h1B65: data = 12'h6FC;
        15'h1B66: data = 12'h706;
        15'h1B67: data = 12'h711;
        15'h1B68: data = 12'h726;
        15'h1B69: data = 12'h734;
        15'h1B6A: data = 12'h734;
        15'h1B6B: data = 12'h744;
        15'h1B6C: data = 12'h751;
        15'h1B6D: data = 12'h75F;
        15'h1B6E: data = 12'h769;
        15'h1B6F: data = 12'h777;
        15'h1B70: data = 12'h77D;
        15'h1B71: data = 12'h790;
        15'h1B72: data = 12'h799;
        15'h1B73: data = 12'h7A0;
        15'h1B74: data = 12'h7A7;
        15'h1B75: data = 12'h7AE;
        15'h1B76: data = 12'h7BC;
        15'h1B77: data = 12'h7C4;
        15'h1B78: data = 12'h7C9;
        15'h1B79: data = 12'h7CE;
        15'h1B7A: data = 12'h7D8;
        15'h1B7B: data = 12'h7DF;
        15'h1B7C: data = 12'h7E9;
        15'h1B7D: data = 12'h7EE;
        15'h1B7E: data = 12'h7F5;
        15'h1B7F: data = 12'h7FD;
        15'h1B80: data = 12'h800;
        15'h1B81: data = 12'h802;
        15'h1B82: data = 12'h80B;
        15'h1B83: data = 12'h80F;
        15'h1B84: data = 12'h81F;
        15'h1B85: data = 12'h08D;
        15'h1B86: data = 12'h095;
        15'h1B87: data = 12'h09B;
        15'h1B88: data = 12'h09B;
        15'h1B89: data = 12'h0A3;
        15'h1B8A: data = 12'h0A3;
        15'h1B8B: data = 12'h0AC;
        15'h1B8C: data = 12'h0AB;
        15'h1B8D: data = 12'h0AD;
        15'h1B8E: data = 12'h0B4;
        15'h1B8F: data = 12'h0B8;
        15'h1B90: data = 12'h0B7;
        15'h1B91: data = 12'h0B7;
        15'h1B92: data = 12'h0BF;
        15'h1B93: data = 12'h0C3;
        15'h1B94: data = 12'h0C8;
        15'h1B95: data = 12'h0C8;
        15'h1B96: data = 12'h0CE;
        15'h1B97: data = 12'h0D0;
        15'h1B98: data = 12'h0D5;
        15'h1B99: data = 12'h0CD;
        15'h1B9A: data = 12'h0CE;
        15'h1B9B: data = 12'h0D0;
        15'h1B9C: data = 12'h0CD;
        15'h1B9D: data = 12'h0CB;
        15'h1B9E: data = 12'h0C0;
        15'h1B9F: data = 12'h0B9;
        15'h1BA0: data = 12'h0AF;
        15'h1BA1: data = 12'h0AD;
        15'h1BA2: data = 12'h0AA;
        15'h1BA3: data = 12'h0A6;
        15'h1BA4: data = 12'h0A5;
        15'h1BA5: data = 12'h0AC;
        15'h1BA6: data = 12'h0A9;
        15'h1BA7: data = 12'h0A5;
        15'h1BA8: data = 12'h0A6;
        15'h1BA9: data = 12'h09E;
        15'h1BAA: data = 12'h094;
        15'h1BAB: data = 12'h089;
        15'h1BAC: data = 12'h07B;
        15'h1BAD: data = 12'h075;
        15'h1BAE: data = 12'h06E;
        15'h1BAF: data = 12'h065;
        15'h1BB0: data = 12'h065;
        15'h1BB1: data = 12'h062;
        15'h1BB2: data = 12'h063;
        15'h1BB3: data = 12'h05B;
        15'h1BB4: data = 12'h051;
        15'h1BB5: data = 12'h03B;
        15'h1BB6: data = 12'h7B9;
        15'h1BB7: data = 12'h7A9;
        15'h1BB8: data = 12'h7A1;
        15'h1BB9: data = 12'h798;
        15'h1BBA: data = 12'h78E;
        15'h1BBB: data = 12'h78D;
        15'h1BBC: data = 12'h780;
        15'h1BBD: data = 12'h776;
        15'h1BBE: data = 12'h761;
        15'h1BBF: data = 12'h753;
        15'h1BC0: data = 12'h73D;
        15'h1BC1: data = 12'h72F;
        15'h1BC2: data = 12'h723;
        15'h1BC3: data = 12'h719;
        15'h1BC4: data = 12'h70F;
        15'h1BC5: data = 12'h70C;
        15'h1BC6: data = 12'h6FF;
        15'h1BC7: data = 12'h6EE;
        15'h1BC8: data = 12'h6E4;
        15'h1BC9: data = 12'h6D1;
        15'h1BCA: data = 12'h6BC;
        15'h1BCB: data = 12'h6AB;
        15'h1BCC: data = 12'h696;
        15'h1BCD: data = 12'h684;
        15'h1BCE: data = 12'h675;
        15'h1BCF: data = 12'h66D;
        15'h1BD0: data = 12'h662;
        15'h1BD1: data = 12'h658;
        15'h1BD2: data = 12'h64B;
        15'h1BD3: data = 12'h639;
        15'h1BD4: data = 12'h62E;
        15'h1BD5: data = 12'h617;
        15'h1BD6: data = 12'h603;
        15'h1BD7: data = 12'h5EC;
        15'h1BD8: data = 12'h5D5;
        15'h1BD9: data = 12'h5BD;
        15'h1BDA: data = 12'h5B2;
        15'h1BDB: data = 12'h5A3;
        15'h1BDC: data = 12'h58E;
        15'h1BDD: data = 12'h581;
        15'h1BDE: data = 12'h56B;
        15'h1BDF: data = 12'h561;
        15'h1BE0: data = 12'h555;
        15'h1BE1: data = 12'h544;
        15'h1BE2: data = 12'h52C;
        15'h1BE3: data = 12'h521;
        15'h1BE4: data = 12'h509;
        15'h1BE5: data = 12'h4F7;
        15'h1BE6: data = 12'h4DE;
        15'h1BE7: data = 12'h4CD;
        15'h1BE8: data = 12'h4B6;
        15'h1BE9: data = 12'h4A3;
        15'h1BEA: data = 12'h487;
        15'h1BEB: data = 12'h470;
        15'h1BEC: data = 12'h454;
        15'h1BED: data = 12'h446;
        15'h1BEE: data = 12'h42F;
        15'h1BEF: data = 12'h417;
        15'h1BF0: data = 12'h3FF;
        15'h1BF1: data = 12'h3E8;
        15'h1BF2: data = 12'h3D4;
        15'h1BF3: data = 12'h3C0;
        15'h1BF4: data = 12'h3AA;
        15'h1BF5: data = 12'h391;
        15'h1BF6: data = 12'h381;
        15'h1BF7: data = 12'h365;
        15'h1BF8: data = 12'h355;
        15'h1BF9: data = 12'h33E;
        15'h1BFA: data = 12'h32B;
        15'h1BFB: data = 12'h31D;
        15'h1BFC: data = 12'h301;
        15'h1BFD: data = 12'h2EA;
        15'h1BFE: data = 12'h2D7;
        15'h1BFF: data = 12'h2C0;
        15'h1C00: data = 12'h2A9;
        15'h1C01: data = 12'h293;
        15'h1C02: data = 12'h280;
        15'h1C03: data = 12'h268;
        15'h1C04: data = 12'h24D;
        15'h1C05: data = 12'h23B;
        15'h1C06: data = 12'h21F;
        15'h1C07: data = 12'h20A;
        15'h1C08: data = 12'h1F4;
        15'h1C09: data = 12'h1DB;
        15'h1C0A: data = 12'h1C2;
        15'h1C0B: data = 12'h1AD;
        15'h1C0C: data = 12'h198;
        15'h1C0D: data = 12'h17E;
        15'h1C0E: data = 12'h169;
        15'h1C0F: data = 12'h151;
        15'h1C10: data = 12'h13C;
        15'h1C11: data = 12'h123;
        15'h1C12: data = 12'h10C;
        15'h1C13: data = 12'h0F3;
        15'h1C14: data = 12'h0DD;
        15'h1C15: data = 12'h0C3;
        15'h1C16: data = 12'h0AC;
        15'h1C17: data = 12'h095;
        15'h1C18: data = 12'h084;
        15'h1C19: data = 12'h064;
        15'h1C1A: data = 12'h050;
        15'h1C1B: data = 12'h52F;
        15'h1C1C: data = 12'h7CE;
        15'h1C1D: data = 12'h7BD;
        15'h1C1E: data = 12'h7A5;
        15'h1C1F: data = 12'h78F;
        15'h1C20: data = 12'h776;
        15'h1C21: data = 12'h75F;
        15'h1C22: data = 12'h74E;
        15'h1C23: data = 12'h737;
        15'h1C24: data = 12'h71D;
        15'h1C25: data = 12'h709;
        15'h1C26: data = 12'h6F1;
        15'h1C27: data = 12'h6DA;
        15'h1C28: data = 12'h6C6;
        15'h1C29: data = 12'h6AD;
        15'h1C2A: data = 12'h698;
        15'h1C2B: data = 12'h684;
        15'h1C2C: data = 12'h66A;
        15'h1C2D: data = 12'h655;
        15'h1C2E: data = 12'h63F;
        15'h1C2F: data = 12'h62D;
        15'h1C30: data = 12'h613;
        15'h1C31: data = 12'h5FB;
        15'h1C32: data = 12'h5E7;
        15'h1C33: data = 12'h5D0;
        15'h1C34: data = 12'h5BF;
        15'h1C35: data = 12'h59E;
        15'h1C36: data = 12'h58A;
        15'h1C37: data = 12'h573;
        15'h1C38: data = 12'h560;
        15'h1C39: data = 12'h54C;
        15'h1C3A: data = 12'h539;
        15'h1C3B: data = 12'h51A;
        15'h1C3C: data = 12'h50B;
        15'h1C3D: data = 12'h4F7;
        15'h1C3E: data = 12'h4DE;
        15'h1C3F: data = 12'h4CC;
        15'h1C40: data = 12'h4B8;
        15'h1C41: data = 12'h4A3;
        15'h1C42: data = 12'h48E;
        15'h1C43: data = 12'h47A;
        15'h1C44: data = 12'h46B;
        15'h1C45: data = 12'h454;
        15'h1C46: data = 12'h447;
        15'h1C47: data = 12'h43B;
        15'h1C48: data = 12'h428;
        15'h1C49: data = 12'h41B;
        15'h1C4A: data = 12'h405;
        15'h1C4B: data = 12'h3FA;
        15'h1C4C: data = 12'h3E8;
        15'h1C4D: data = 12'h3D3;
        15'h1C4E: data = 12'h3C4;
        15'h1C4F: data = 12'h3B1;
        15'h1C50: data = 12'h39E;
        15'h1C51: data = 12'h390;
        15'h1C52: data = 12'h379;
        15'h1C53: data = 12'h36A;
        15'h1C54: data = 12'h359;
        15'h1C55: data = 12'h344;
        15'h1C56: data = 12'h332;
        15'h1C57: data = 12'h31D;
        15'h1C58: data = 12'h30F;
        15'h1C59: data = 12'h2FD;
        15'h1C5A: data = 12'h2EE;
        15'h1C5B: data = 12'h2E3;
        15'h1C5C: data = 12'h2D4;
        15'h1C5D: data = 12'h2CE;
        15'h1C5E: data = 12'h2C2;
        15'h1C5F: data = 12'h2B6;
        15'h1C60: data = 12'h2A8;
        15'h1C61: data = 12'h2A2;
        15'h1C62: data = 12'h295;
        15'h1C63: data = 12'h283;
        15'h1C64: data = 12'h27D;
        15'h1C65: data = 12'h26D;
        15'h1C66: data = 12'h261;
        15'h1C67: data = 12'h24C;
        15'h1C68: data = 12'h244;
        15'h1C69: data = 12'h230;
        15'h1C6A: data = 12'h223;
        15'h1C6B: data = 12'h215;
        15'h1C6C: data = 12'h212;
        15'h1C6D: data = 12'h208;
        15'h1C6E: data = 12'h201;
        15'h1C6F: data = 12'h1F4;
        15'h1C70: data = 12'h1F4;
        15'h1C71: data = 12'h1EE;
        15'h1C72: data = 12'h1E9;
        15'h1C73: data = 12'h1E1;
        15'h1C74: data = 12'h1D5;
        15'h1C75: data = 12'h1CE;
        15'h1C76: data = 12'h1C4;
        15'h1C77: data = 12'h1BF;
        15'h1C78: data = 12'h1B4;
        15'h1C79: data = 12'h1A7;
        15'h1C7A: data = 12'h19C;
        15'h1C7B: data = 12'h192;
        15'h1C7C: data = 12'h195;
        15'h1C7D: data = 12'h18E;
        15'h1C7E: data = 12'h187;
        15'h1C7F: data = 12'h187;
        15'h1C80: data = 12'h188;
        15'h1C81: data = 12'h183;
        15'h1C82: data = 12'h185;
        15'h1C83: data = 12'h17F;
        15'h1C84: data = 12'h180;
        15'h1C85: data = 12'h178;
        15'h1C86: data = 12'h176;
        15'h1C87: data = 12'h174;
        15'h1C88: data = 12'h164;
        15'h1C89: data = 12'h162;
        15'h1C8A: data = 12'h15E;
        15'h1C8B: data = 12'h15C;
        15'h1C8C: data = 12'h154;
        15'h1C8D: data = 12'h157;
        15'h1C8E: data = 12'h158;
        15'h1C8F: data = 12'h15D;
        15'h1C90: data = 12'h161;
        15'h1C91: data = 12'h164;
        15'h1C92: data = 12'h168;
        15'h1C93: data = 12'h172;
        15'h1C94: data = 12'h16D;
        15'h1C95: data = 12'h16E;
        15'h1C96: data = 12'h16B;
        15'h1C97: data = 12'h169;
        15'h1C98: data = 12'h16B;
        15'h1C99: data = 12'h168;
        15'h1C9A: data = 12'h16B;
        15'h1C9B: data = 12'h16E;
        15'h1C9C: data = 12'h16C;
        15'h1C9D: data = 12'h176;
        15'h1C9E: data = 12'h17B;
        15'h1C9F: data = 12'h182;
        15'h1CA0: data = 12'h18A;
        15'h1CA1: data = 12'h18F;
        15'h1CA2: data = 12'h19D;
        15'h1CA3: data = 12'h1A3;
        15'h1CA4: data = 12'h1AC;
        15'h1CA5: data = 12'h1B3;
        15'h1CA6: data = 12'h1B3;
        15'h1CA7: data = 12'h1B7;
        15'h1CA8: data = 12'h1BE;
        15'h1CA9: data = 12'h1C2;
        15'h1CAA: data = 12'h1C5;
        15'h1CAB: data = 12'h1CC;
        15'h1CAC: data = 12'h1D0;
        15'h1CAD: data = 12'h1D7;
        15'h1CAE: data = 12'h1E2;
        15'h1CAF: data = 12'h1ED;
        15'h1CB0: data = 12'h1FB;
        15'h1CB1: data = 12'h207;
        15'h1CB2: data = 12'h217;
        15'h1CB3: data = 12'h21D;
        15'h1CB4: data = 12'h22F;
        15'h1CB5: data = 12'h238;
        15'h1CB6: data = 12'h245;
        15'h1CB7: data = 12'h24C;
        15'h1CB8: data = 12'h25C;
        15'h1CB9: data = 12'h262;
        15'h1CBA: data = 12'h26E;
        15'h1CBB: data = 12'h274;
        15'h1CBC: data = 12'h27F;
        15'h1CBD: data = 12'h287;
        15'h1CBE: data = 12'h292;
        15'h1CBF: data = 12'h2A3;
        15'h1CC0: data = 12'h2AE;
        15'h1CC1: data = 12'h2BD;
        15'h1CC2: data = 12'h2D1;
        15'h1CC3: data = 12'h2DE;
        15'h1CC4: data = 12'h2F1;
        15'h1CC5: data = 12'h304;
        15'h1CC6: data = 12'h31A;
        15'h1CC7: data = 12'h329;
        15'h1CC8: data = 12'h337;
        15'h1CC9: data = 12'h347;
        15'h1CCA: data = 12'h355;
        15'h1CCB: data = 12'h366;
        15'h1CCC: data = 12'h373;
        15'h1CCD: data = 12'h381;
        15'h1CCE: data = 12'h394;
        15'h1CCF: data = 12'h39B;
        15'h1CD0: data = 12'h3AD;
        15'h1CD1: data = 12'h3BB;
        15'h1CD2: data = 12'h3C8;
        15'h1CD3: data = 12'h3DF;
        15'h1CD4: data = 12'h3EE;
        15'h1CD5: data = 12'h3FE;
        15'h1CD6: data = 12'h414;
        15'h1CD7: data = 12'h426;
        15'h1CD8: data = 12'h43C;
        15'h1CD9: data = 12'h451;
        15'h1CDA: data = 12'h466;
        15'h1CDB: data = 12'h47E;
        15'h1CDC: data = 12'h492;
        15'h1CDD: data = 12'h4AB;
        15'h1CDE: data = 12'h4BC;
        15'h1CDF: data = 12'h4CE;
        15'h1CE0: data = 12'h4E5;
        15'h1CE1: data = 12'h4F6;
        15'h1CE2: data = 12'h50B;
        15'h1CE3: data = 12'h51A;
        15'h1CE4: data = 12'h52C;
        15'h1CE5: data = 12'h541;
        15'h1CE6: data = 12'h554;
        15'h1CE7: data = 12'h561;
        15'h1CE8: data = 12'h575;
        15'h1CE9: data = 12'h58B;
        15'h1CEA: data = 12'h5A0;
        15'h1CEB: data = 12'h5B7;
        15'h1CEC: data = 12'h5CB;
        15'h1CED: data = 12'h5E3;
        15'h1CEE: data = 12'h5FB;
        15'h1CEF: data = 12'h61A;
        15'h1CF0: data = 12'h630;
        15'h1CF1: data = 12'h645;
        15'h1CF2: data = 12'h65F;
        15'h1CF3: data = 12'h675;
        15'h1CF4: data = 12'h693;
        15'h1CF5: data = 12'h6A5;
        15'h1CF6: data = 12'h6BB;
        15'h1CF7: data = 12'h6CE;
        15'h1CF8: data = 12'h6E3;
        15'h1CF9: data = 12'h6F8;
        15'h1CFA: data = 12'h70F;
        15'h1CFB: data = 12'h724;
        15'h1CFC: data = 12'h737;
        15'h1CFD: data = 12'h747;
        15'h1CFE: data = 12'h75E;
        15'h1CFF: data = 12'h775;
        15'h1D00: data = 12'h78D;
        15'h1D01: data = 12'h79F;
        15'h1D02: data = 12'h7B8;
        15'h1D03: data = 12'h7D0;
        15'h1D04: data = 12'h7E7;
        15'h1D05: data = 12'h7FD;
        15'h1D06: data = 12'h104;
        15'h1D07: data = 12'h089;
        15'h1D08: data = 12'h09F;
        15'h1D09: data = 12'h0B1;
        15'h1D0A: data = 12'h0D0;
        15'h1D0B: data = 12'h0E9;
        15'h1D0C: data = 12'h101;
        15'h1D0D: data = 12'h112;
        15'h1D0E: data = 12'h129;
        15'h1D0F: data = 12'h140;
        15'h1D10: data = 12'h158;
        15'h1D11: data = 12'h16F;
        15'h1D12: data = 12'h180;
        15'h1D13: data = 12'h19B;
        15'h1D14: data = 12'h1B1;
        15'h1D15: data = 12'h1BF;
        15'h1D16: data = 12'h1D7;
        15'h1D17: data = 12'h1F1;
        15'h1D18: data = 12'h207;
        15'h1D19: data = 12'h219;
        15'h1D1A: data = 12'h231;
        15'h1D1B: data = 12'h249;
        15'h1D1C: data = 12'h25F;
        15'h1D1D: data = 12'h276;
        15'h1D1E: data = 12'h28C;
        15'h1D1F: data = 12'h2A2;
        15'h1D20: data = 12'h2C0;
        15'h1D21: data = 12'h2D6;
        15'h1D22: data = 12'h2F1;
        15'h1D23: data = 12'h304;
        15'h1D24: data = 12'h322;
        15'h1D25: data = 12'h32E;
        15'h1D26: data = 12'h34A;
        15'h1D27: data = 12'h364;
        15'h1D28: data = 12'h37E;
        15'h1D29: data = 12'h396;
        15'h1D2A: data = 12'h3AA;
        15'h1D2B: data = 12'h3C3;
        15'h1D2C: data = 12'h3DB;
        15'h1D2D: data = 12'h3EF;
        15'h1D2E: data = 12'h3FF;
        15'h1D2F: data = 12'h417;
        15'h1D30: data = 12'h42E;
        15'h1D31: data = 12'h442;
        15'h1D32: data = 12'h456;
        15'h1D33: data = 12'h468;
        15'h1D34: data = 12'h480;
        15'h1D35: data = 12'h497;
        15'h1D36: data = 12'h4A9;
        15'h1D37: data = 12'h4BC;
        15'h1D38: data = 12'h4C8;
        15'h1D39: data = 12'h4E0;
        15'h1D3A: data = 12'h4F5;
        15'h1D3B: data = 12'h508;
        15'h1D3C: data = 12'h514;
        15'h1D3D: data = 12'h529;
        15'h1D3E: data = 12'h53B;
        15'h1D3F: data = 12'h548;
        15'h1D40: data = 12'h55E;
        15'h1D41: data = 12'h56C;
        15'h1D42: data = 12'h581;
        15'h1D43: data = 12'h596;
        15'h1D44: data = 12'h5A3;
        15'h1D45: data = 12'h5B7;
        15'h1D46: data = 12'h5C5;
        15'h1D47: data = 12'h5D6;
        15'h1D48: data = 12'h5F0;
        15'h1D49: data = 12'h5FD;
        15'h1D4A: data = 12'h60A;
        15'h1D4B: data = 12'h619;
        15'h1D4C: data = 12'h62A;
        15'h1D4D: data = 12'h638;
        15'h1D4E: data = 12'h64E;
        15'h1D4F: data = 12'h660;
        15'h1D50: data = 12'h672;
        15'h1D51: data = 12'h67F;
        15'h1D52: data = 12'h692;
        15'h1D53: data = 12'h6A0;
        15'h1D54: data = 12'h6AE;
        15'h1D55: data = 12'h6C1;
        15'h1D56: data = 12'h6CC;
        15'h1D57: data = 12'h6D8;
        15'h1D58: data = 12'h6EA;
        15'h1D59: data = 12'h6FA;
        15'h1D5A: data = 12'h705;
        15'h1D5B: data = 12'h714;
        15'h1D5C: data = 12'h725;
        15'h1D5D: data = 12'h731;
        15'h1D5E: data = 12'h737;
        15'h1D5F: data = 12'h741;
        15'h1D60: data = 12'h751;
        15'h1D61: data = 12'h762;
        15'h1D62: data = 12'h769;
        15'h1D63: data = 12'h776;
        15'h1D64: data = 12'h77F;
        15'h1D65: data = 12'h78C;
        15'h1D66: data = 12'h794;
        15'h1D67: data = 12'h79B;
        15'h1D68: data = 12'h7A2;
        15'h1D69: data = 12'h7B1;
        15'h1D6A: data = 12'h7B8;
        15'h1D6B: data = 12'h7C0;
        15'h1D6C: data = 12'h7C9;
        15'h1D6D: data = 12'h7CD;
        15'h1D6E: data = 12'h7D4;
        15'h1D6F: data = 12'h7DF;
        15'h1D70: data = 12'h7E5;
        15'h1D71: data = 12'h7ED;
        15'h1D72: data = 12'h7F7;
        15'h1D73: data = 12'h7F9;
        15'h1D74: data = 12'h801;
        15'h1D75: data = 12'h801;
        15'h1D76: data = 12'h803;
        15'h1D77: data = 12'h80D;
        15'h1D78: data = 12'h885;
        15'h1D79: data = 12'h08A;
        15'h1D7A: data = 12'h098;
        15'h1D7B: data = 12'h09B;
        15'h1D7C: data = 12'h09B;
        15'h1D7D: data = 12'h0A2;
        15'h1D7E: data = 12'h0A6;
        15'h1D7F: data = 12'h0AC;
        15'h1D80: data = 12'h0AB;
        15'h1D81: data = 12'h0AA;
        15'h1D82: data = 12'h0B2;
        15'h1D83: data = 12'h0B5;
        15'h1D84: data = 12'h0B7;
        15'h1D85: data = 12'h0BA;
        15'h1D86: data = 12'h0C2;
        15'h1D87: data = 12'h0C3;
        15'h1D88: data = 12'h0C5;
        15'h1D89: data = 12'h0CC;
        15'h1D8A: data = 12'h0CD;
        15'h1D8B: data = 12'h0D2;
        15'h1D8C: data = 12'h0D1;
        15'h1D8D: data = 12'h0CC;
        15'h1D8E: data = 12'h0CE;
        15'h1D8F: data = 12'h0CC;
        15'h1D90: data = 12'h0CB;
        15'h1D91: data = 12'h0C9;
        15'h1D92: data = 12'h0BD;
        15'h1D93: data = 12'h0BC;
        15'h1D94: data = 12'h0B1;
        15'h1D95: data = 12'h0AC;
        15'h1D96: data = 12'h0A9;
        15'h1D97: data = 12'h0A8;
        15'h1D98: data = 12'h0A3;
        15'h1D99: data = 12'h0AC;
        15'h1D9A: data = 12'h0AA;
        15'h1D9B: data = 12'h0A4;
        15'h1D9C: data = 12'h0A5;
        15'h1D9D: data = 12'h09F;
        15'h1D9E: data = 12'h096;
        15'h1D9F: data = 12'h08A;
        15'h1DA0: data = 12'h079;
        15'h1DA1: data = 12'h077;
        15'h1DA2: data = 12'h06A;
        15'h1DA3: data = 12'h065;
        15'h1DA4: data = 12'h064;
        15'h1DA5: data = 12'h064;
        15'h1DA6: data = 12'h062;
        15'h1DA7: data = 12'h05A;
        15'h1DA8: data = 12'h04E;
        15'h1DA9: data = 12'h040;
        15'h1DAA: data = 12'h7BB;
        15'h1DAB: data = 12'h7A9;
        15'h1DAC: data = 12'h7A2;
        15'h1DAD: data = 12'h793;
        15'h1DAE: data = 12'h78F;
        15'h1DAF: data = 12'h78E;
        15'h1DB0: data = 12'h77F;
        15'h1DB1: data = 12'h773;
        15'h1DB2: data = 12'h75F;
        15'h1DB3: data = 12'h750;
        15'h1DB4: data = 12'h73A;
        15'h1DB5: data = 12'h72C;
        15'h1DB6: data = 12'h723;
        15'h1DB7: data = 12'h714;
        15'h1DB8: data = 12'h70C;
        15'h1DB9: data = 12'h70A;
        15'h1DBA: data = 12'h6FD;
        15'h1DBB: data = 12'h6EF;
        15'h1DBC: data = 12'h6E4;
        15'h1DBD: data = 12'h6CD;
        15'h1DBE: data = 12'h6B7;
        15'h1DBF: data = 12'h6A7;
        15'h1DC0: data = 12'h696;
        15'h1DC1: data = 12'h687;
        15'h1DC2: data = 12'h67D;
        15'h1DC3: data = 12'h66E;
        15'h1DC4: data = 12'h662;
        15'h1DC5: data = 12'h656;
        15'h1DC6: data = 12'h649;
        15'h1DC7: data = 12'h638;
        15'h1DC8: data = 12'h630;
        15'h1DC9: data = 12'h615;
        15'h1DCA: data = 12'h600;
        15'h1DCB: data = 12'h5ED;
        15'h1DCC: data = 12'h5D2;
        15'h1DCD: data = 12'h5BE;
        15'h1DCE: data = 12'h5AD;
        15'h1DCF: data = 12'h5A0;
        15'h1DD0: data = 12'h58E;
        15'h1DD1: data = 12'h580;
        15'h1DD2: data = 12'h571;
        15'h1DD3: data = 12'h564;
        15'h1DD4: data = 12'h555;
        15'h1DD5: data = 12'h546;
        15'h1DD6: data = 12'h52E;
        15'h1DD7: data = 12'h51D;
        15'h1DD8: data = 12'h50A;
        15'h1DD9: data = 12'h4F7;
        15'h1DDA: data = 12'h4DB;
        15'h1DDB: data = 12'h4C8;
        15'h1DDC: data = 12'h4B5;
        15'h1DDD: data = 12'h49D;
        15'h1DDE: data = 12'h485;
        15'h1DDF: data = 12'h46E;
        15'h1DE0: data = 12'h457;
        15'h1DE1: data = 12'h444;
        15'h1DE2: data = 12'h42B;
        15'h1DE3: data = 12'h416;
        15'h1DE4: data = 12'h3FE;
        15'h1DE5: data = 12'h3E5;
        15'h1DE6: data = 12'h3D6;
        15'h1DE7: data = 12'h3C2;
        15'h1DE8: data = 12'h3AD;
        15'h1DE9: data = 12'h395;
        15'h1DEA: data = 12'h37F;
        15'h1DEB: data = 12'h369;
        15'h1DEC: data = 12'h357;
        15'h1DED: data = 12'h342;
        15'h1DEE: data = 12'h32D;
        15'h1DEF: data = 12'h31B;
        15'h1DF0: data = 12'h300;
        15'h1DF1: data = 12'h2ED;
        15'h1DF2: data = 12'h2D6;
        15'h1DF3: data = 12'h2C2;
        15'h1DF4: data = 12'h2A8;
        15'h1DF5: data = 12'h291;
        15'h1DF6: data = 12'h27D;
        15'h1DF7: data = 12'h26A;
        15'h1DF8: data = 12'h24D;
        15'h1DF9: data = 12'h23A;
        15'h1DFA: data = 12'h21D;
        15'h1DFB: data = 12'h209;
        15'h1DFC: data = 12'h1F6;
        15'h1DFD: data = 12'h1DD;
        15'h1DFE: data = 12'h1C1;
        15'h1DFF: data = 12'h1AC;
        15'h1E00: data = 12'h197;
        15'h1E01: data = 12'h180;
        15'h1E02: data = 12'h168;
        15'h1E03: data = 12'h152;
        15'h1E04: data = 12'h13C;
        15'h1E05: data = 12'h120;
        15'h1E06: data = 12'h109;
        15'h1E07: data = 12'h0F5;
        15'h1E08: data = 12'h0DD;
        15'h1E09: data = 12'h0C4;
        15'h1E0A: data = 12'h0A8;
        15'h1E0B: data = 12'h095;
        15'h1E0C: data = 12'h081;
        15'h1E0D: data = 12'h066;
        15'h1E0E: data = 12'h052;
        15'h1E0F: data = 12'h4C6;
        15'h1E10: data = 12'h7CF;
        15'h1E11: data = 12'h7BF;
        15'h1E12: data = 12'h7A6;
        15'h1E13: data = 12'h78E;
        15'h1E14: data = 12'h779;
        15'h1E15: data = 12'h760;
        15'h1E16: data = 12'h74C;
        15'h1E17: data = 12'h736;
        15'h1E18: data = 12'h71E;
        15'h1E19: data = 12'h709;
        15'h1E1A: data = 12'h6F1;
        15'h1E1B: data = 12'h6DB;
        15'h1E1C: data = 12'h6C4;
        15'h1E1D: data = 12'h6B1;
        15'h1E1E: data = 12'h694;
        15'h1E1F: data = 12'h683;
        15'h1E20: data = 12'h66D;
        15'h1E21: data = 12'h658;
        15'h1E22: data = 12'h63F;
        15'h1E23: data = 12'h62C;
        15'h1E24: data = 12'h614;
        15'h1E25: data = 12'h5FE;
        15'h1E26: data = 12'h5E6;
        15'h1E27: data = 12'h5CE;
        15'h1E28: data = 12'h5BD;
        15'h1E29: data = 12'h59F;
        15'h1E2A: data = 12'h589;
        15'h1E2B: data = 12'h576;
        15'h1E2C: data = 12'h565;
        15'h1E2D: data = 12'h54F;
        15'h1E2E: data = 12'h536;
        15'h1E2F: data = 12'h51A;
        15'h1E30: data = 12'h50E;
        15'h1E31: data = 12'h4F5;
        15'h1E32: data = 12'h4DE;
        15'h1E33: data = 12'h4CD;
        15'h1E34: data = 12'h4B8;
        15'h1E35: data = 12'h4A5;
        15'h1E36: data = 12'h48F;
        15'h1E37: data = 12'h47D;
        15'h1E38: data = 12'h46A;
        15'h1E39: data = 12'h458;
        15'h1E3A: data = 12'h44A;
        15'h1E3B: data = 12'h43E;
        15'h1E3C: data = 12'h429;
        15'h1E3D: data = 12'h418;
        15'h1E3E: data = 12'h409;
        15'h1E3F: data = 12'h3F8;
        15'h1E40: data = 12'h3EA;
        15'h1E41: data = 12'h3D4;
        15'h1E42: data = 12'h3C0;
        15'h1E43: data = 12'h3B2;
        15'h1E44: data = 12'h39F;
        15'h1E45: data = 12'h392;
        15'h1E46: data = 12'h37E;
        15'h1E47: data = 12'h366;
        15'h1E48: data = 12'h359;
        15'h1E49: data = 12'h345;
        15'h1E4A: data = 12'h32E;
        15'h1E4B: data = 12'h31F;
        15'h1E4C: data = 12'h311;
        15'h1E4D: data = 12'h2FB;
        15'h1E4E: data = 12'h2F0;
        15'h1E4F: data = 12'h2DF;
        15'h1E50: data = 12'h2D3;
        15'h1E51: data = 12'h2D0;
        15'h1E52: data = 12'h2C7;
        15'h1E53: data = 12'h2B7;
        15'h1E54: data = 12'h2AB;
        15'h1E55: data = 12'h2A1;
        15'h1E56: data = 12'h295;
        15'h1E57: data = 12'h287;
        15'h1E58: data = 12'h27C;
        15'h1E59: data = 12'h26C;
        15'h1E5A: data = 12'h264;
        15'h1E5B: data = 12'h250;
        15'h1E5C: data = 12'h243;
        15'h1E5D: data = 12'h22F;
        15'h1E5E: data = 12'h226;
        15'h1E5F: data = 12'h216;
        15'h1E60: data = 12'h211;
        15'h1E61: data = 12'h206;
        15'h1E62: data = 12'h201;
        15'h1E63: data = 12'h1F8;
        15'h1E64: data = 12'h1F3;
        15'h1E65: data = 12'h1EF;
        15'h1E66: data = 12'h1EC;
        15'h1E67: data = 12'h1E6;
        15'h1E68: data = 12'h1D7;
        15'h1E69: data = 12'h1CE;
        15'h1E6A: data = 12'h1C5;
        15'h1E6B: data = 12'h1C1;
        15'h1E6C: data = 12'h1B6;
        15'h1E6D: data = 12'h1AA;
        15'h1E6E: data = 12'h19D;
        15'h1E6F: data = 12'h195;
        15'h1E70: data = 12'h192;
        15'h1E71: data = 12'h18B;
        15'h1E72: data = 12'h186;
        15'h1E73: data = 12'h185;
        15'h1E74: data = 12'h188;
        15'h1E75: data = 12'h184;
        15'h1E76: data = 12'h184;
        15'h1E77: data = 12'h181;
        15'h1E78: data = 12'h181;
        15'h1E79: data = 12'h177;
        15'h1E7A: data = 12'h175;
        15'h1E7B: data = 12'h175;
        15'h1E7C: data = 12'h168;
        15'h1E7D: data = 12'h163;
        15'h1E7E: data = 12'h15F;
        15'h1E7F: data = 12'h15E;
        15'h1E80: data = 12'h153;
        15'h1E81: data = 12'h157;
        15'h1E82: data = 12'h159;
        15'h1E83: data = 12'h15A;
        15'h1E84: data = 12'h161;
        15'h1E85: data = 12'h163;
        15'h1E86: data = 12'h16A;
        15'h1E87: data = 12'h16F;
        15'h1E88: data = 12'h173;
        15'h1E89: data = 12'h16F;
        15'h1E8A: data = 12'h16C;
        15'h1E8B: data = 12'h16B;
        15'h1E8C: data = 12'h171;
        15'h1E8D: data = 12'h167;
        15'h1E8E: data = 12'h169;
        15'h1E8F: data = 12'h16B;
        15'h1E90: data = 12'h16B;
        15'h1E91: data = 12'h175;
        15'h1E92: data = 12'h17D;
        15'h1E93: data = 12'h183;
        15'h1E94: data = 12'h18C;
        15'h1E95: data = 12'h191;
        15'h1E96: data = 12'h19D;
        15'h1E97: data = 12'h1A8;
        15'h1E98: data = 12'h1AD;
        15'h1E99: data = 12'h1B0;
        15'h1E9A: data = 12'h1B3;
        15'h1E9B: data = 12'h1BA;
        15'h1E9C: data = 12'h1BF;
        15'h1E9D: data = 12'h1C3;
        15'h1E9E: data = 12'h1C7;
        15'h1E9F: data = 12'h1CB;
        15'h1EA0: data = 12'h1D2;
        15'h1EA1: data = 12'h1DA;
        15'h1EA2: data = 12'h1E1;
        15'h1EA3: data = 12'h1EE;
        15'h1EA4: data = 12'h1FA;
        15'h1EA5: data = 12'h205;
        15'h1EA6: data = 12'h218;
        15'h1EA7: data = 12'h21E;
        15'h1EA8: data = 12'h22F;
        15'h1EA9: data = 12'h23A;
        15'h1EAA: data = 12'h247;
        15'h1EAB: data = 12'h24C;
        15'h1EAC: data = 12'h25C;
        15'h1EAD: data = 12'h264;
        15'h1EAE: data = 12'h271;
        15'h1EAF: data = 12'h273;
        15'h1EB0: data = 12'h280;
        15'h1EB1: data = 12'h286;
        15'h1EB2: data = 12'h291;
        15'h1EB3: data = 12'h2A3;
        15'h1EB4: data = 12'h2AF;
        15'h1EB5: data = 12'h2BF;
        15'h1EB6: data = 12'h2D0;
        15'h1EB7: data = 12'h2DF;
        15'h1EB8: data = 12'h2F0;
        15'h1EB9: data = 12'h301;
        15'h1EBA: data = 12'h316;
        15'h1EBB: data = 12'h328;
        15'h1EBC: data = 12'h338;
        15'h1EBD: data = 12'h346;
        15'h1EBE: data = 12'h357;
        15'h1EBF: data = 12'h365;
        15'h1EC0: data = 12'h374;
        15'h1EC1: data = 12'h383;
        15'h1EC2: data = 12'h397;
        15'h1EC3: data = 12'h399;
        15'h1EC4: data = 12'h3B0;
        15'h1EC5: data = 12'h3B9;
        15'h1EC6: data = 12'h3C9;
        15'h1EC7: data = 12'h3DD;
        15'h1EC8: data = 12'h3EE;
        15'h1EC9: data = 12'h3FB;
        15'h1ECA: data = 12'h413;
        15'h1ECB: data = 12'h428;
        15'h1ECC: data = 12'h43D;
        15'h1ECD: data = 12'h453;
        15'h1ECE: data = 12'h467;
        15'h1ECF: data = 12'h480;
        15'h1ED0: data = 12'h492;
        15'h1ED1: data = 12'h4AB;
        15'h1ED2: data = 12'h4B9;
        15'h1ED3: data = 12'h4D2;
        15'h1ED4: data = 12'h4E3;
        15'h1ED5: data = 12'h4F5;
        15'h1ED6: data = 12'h509;
        15'h1ED7: data = 12'h51B;
        15'h1ED8: data = 12'h52A;
        15'h1ED9: data = 12'h53F;
        15'h1EDA: data = 12'h553;
        15'h1EDB: data = 12'h566;
        15'h1EDC: data = 12'h574;
        15'h1EDD: data = 12'h58C;
        15'h1EDE: data = 12'h5A0;
        15'h1EDF: data = 12'h5B7;
        15'h1EE0: data = 12'h5CC;
        15'h1EE1: data = 12'h5E1;
        15'h1EE2: data = 12'h5FB;
        15'h1EE3: data = 12'h616;
        15'h1EE4: data = 12'h62D;
        15'h1EE5: data = 12'h643;
        15'h1EE6: data = 12'h660;
        15'h1EE7: data = 12'h677;
        15'h1EE8: data = 12'h690;
        15'h1EE9: data = 12'h6A1;
        15'h1EEA: data = 12'h6BB;
        15'h1EEB: data = 12'h6D2;
        15'h1EEC: data = 12'h6E1;
        15'h1EED: data = 12'h6F6;
        15'h1EEE: data = 12'h70D;
        15'h1EEF: data = 12'h724;
        15'h1EF0: data = 12'h73A;
        15'h1EF1: data = 12'h74B;
        15'h1EF2: data = 12'h75D;
        15'h1EF3: data = 12'h773;
        15'h1EF4: data = 12'h78D;
        15'h1EF5: data = 12'h7A0;
        15'h1EF6: data = 12'h7B8;
        15'h1EF7: data = 12'h7D2;
        15'h1EF8: data = 12'h7E6;
        15'h1EF9: data = 12'h800;
        15'h1EFA: data = 12'h06C;
        15'h1EFB: data = 12'h088;
        15'h1EFC: data = 12'h0A0;
        15'h1EFD: data = 12'h0B3;
        15'h1EFE: data = 12'h0D1;
        15'h1EFF: data = 12'h0E9;
        15'h1F00: data = 12'h100;
        15'h1F01: data = 12'h111;
        15'h1F02: data = 12'h12E;
        15'h1F03: data = 12'h144;
        15'h1F04: data = 12'h158;
        15'h1F05: data = 12'h16D;
        15'h1F06: data = 12'h181;
        15'h1F07: data = 12'h19D;
        15'h1F08: data = 12'h1B5;
        15'h1F09: data = 12'h1C0;
        15'h1F0A: data = 12'h1DC;
        15'h1F0B: data = 12'h1F0;
        15'h1F0C: data = 12'h205;
        15'h1F0D: data = 12'h218;
        15'h1F0E: data = 12'h232;
        15'h1F0F: data = 12'h249;
        15'h1F10: data = 12'h25D;
        15'h1F11: data = 12'h277;
        15'h1F12: data = 12'h289;
        15'h1F13: data = 12'h2A7;
        15'h1F14: data = 12'h2BF;
        15'h1F15: data = 12'h2D1;
        15'h1F16: data = 12'h2EF;
        15'h1F17: data = 12'h305;
        15'h1F18: data = 12'h320;
        15'h1F19: data = 12'h332;
        15'h1F1A: data = 12'h34A;
        15'h1F1B: data = 12'h366;
        15'h1F1C: data = 12'h37C;
        15'h1F1D: data = 12'h398;
        15'h1F1E: data = 12'h3AB;
        15'h1F1F: data = 12'h3C3;
        15'h1F20: data = 12'h3DD;
        15'h1F21: data = 12'h3F0;
        15'h1F22: data = 12'h402;
        15'h1F23: data = 12'h417;
        15'h1F24: data = 12'h42F;
        15'h1F25: data = 12'h445;
        15'h1F26: data = 12'h454;
        15'h1F27: data = 12'h46A;
        15'h1F28: data = 12'h47E;
        15'h1F29: data = 12'h498;
        15'h1F2A: data = 12'h4A8;
        15'h1F2B: data = 12'h4BC;
        15'h1F2C: data = 12'h4CC;
        15'h1F2D: data = 12'h4DC;
        15'h1F2E: data = 12'h4F0;
        15'h1F2F: data = 12'h505;
        15'h1F30: data = 12'h510;
        15'h1F31: data = 12'h526;
        15'h1F32: data = 12'h53C;
        15'h1F33: data = 12'h547;
        15'h1F34: data = 12'h55E;
        15'h1F35: data = 12'h56B;
        15'h1F36: data = 12'h582;
        15'h1F37: data = 12'h591;
        15'h1F38: data = 12'h5A4;
        15'h1F39: data = 12'h5BA;
        15'h1F3A: data = 12'h5C4;
        15'h1F3B: data = 12'h5D4;
        15'h1F3C: data = 12'h5E9;
        15'h1F3D: data = 12'h5FB;
        15'h1F3E: data = 12'h60D;
        15'h1F3F: data = 12'h61D;
        15'h1F40: data = 12'h62B;
        15'h1F41: data = 12'h63B;
        15'h1F42: data = 12'h64E;
        15'h1F43: data = 12'h661;
        15'h1F44: data = 12'h671;
        15'h1F45: data = 12'h680;
        15'h1F46: data = 12'h693;
        15'h1F47: data = 12'h6A1;
        15'h1F48: data = 12'h6AF;
        15'h1F49: data = 12'h6C0;
        15'h1F4A: data = 12'h6D1;
        15'h1F4B: data = 12'h6DD;
        15'h1F4C: data = 12'h6EA;
        15'h1F4D: data = 12'h6F9;
        15'h1F4E: data = 12'h702;
        15'h1F4F: data = 12'h715;
        15'h1F50: data = 12'h725;
        15'h1F51: data = 12'h734;
        15'h1F52: data = 12'h737;
        15'h1F53: data = 12'h744;
        15'h1F54: data = 12'h74E;
        15'h1F55: data = 12'h75F;
        15'h1F56: data = 12'h768;
        15'h1F57: data = 12'h778;
        15'h1F58: data = 12'h77D;
        15'h1F59: data = 12'h78E;
        15'h1F5A: data = 12'h795;
        15'h1F5B: data = 12'h79D;
        15'h1F5C: data = 12'h7A5;
        15'h1F5D: data = 12'h7B2;
        15'h1F5E: data = 12'h7BB;
        15'h1F5F: data = 12'h7C2;
        15'h1F60: data = 12'h7C7;
        15'h1F61: data = 12'h7D0;
        15'h1F62: data = 12'h7DA;
        15'h1F63: data = 12'h7DD;
        15'h1F64: data = 12'h7E4;
        15'h1F65: data = 12'h7EF;
        15'h1F66: data = 12'h7F4;
        15'h1F67: data = 12'h7FD;
        15'h1F68: data = 12'h800;
        15'h1F69: data = 12'h802;
        15'h1F6A: data = 12'h809;
        15'h1F6B: data = 12'h073;
        15'h1F6C: data = 12'h08F;
        15'h1F6D: data = 12'h090;
        15'h1F6E: data = 12'h09A;
        15'h1F6F: data = 12'h09D;
        15'h1F70: data = 12'h09B;
        15'h1F71: data = 12'h0A3;
        15'h1F72: data = 12'h0A6;
        15'h1F73: data = 12'h0B0;
        15'h1F74: data = 12'h0B1;
        15'h1F75: data = 12'h0AC;
        15'h1F76: data = 12'h0B8;
        15'h1F77: data = 12'h0B8;
        15'h1F78: data = 12'h0BD;
        15'h1F79: data = 12'h0BA;
        15'h1F7A: data = 12'h0C6;
        15'h1F7B: data = 12'h0C9;
        15'h1F7C: data = 12'h0CF;
        15'h1F7D: data = 12'h0D2;
        15'h1F7E: data = 12'h0D2;
        15'h1F7F: data = 12'h0D8;
        15'h1F80: data = 12'h0D7;
        15'h1F81: data = 12'h0CD;
        15'h1F82: data = 12'h0CC;
        15'h1F83: data = 12'h0CB;
        15'h1F84: data = 12'h0C8;
        15'h1F85: data = 12'h0C5;
        15'h1F86: data = 12'h0BC;
        15'h1F87: data = 12'h0B6;
        15'h1F88: data = 12'h0AC;
        15'h1F89: data = 12'h0AC;
        15'h1F8A: data = 12'h0A9;
        15'h1F8B: data = 12'h0AB;
        15'h1F8C: data = 12'h0AF;
        15'h1F8D: data = 12'h0B3;
        15'h1F8E: data = 12'h0AD;
        15'h1F8F: data = 12'h0A5;
        15'h1F90: data = 12'h0A5;
        15'h1F91: data = 12'h099;
        15'h1F92: data = 12'h090;
        15'h1F93: data = 12'h080;
        15'h1F94: data = 12'h075;
        15'h1F95: data = 12'h075;
        15'h1F96: data = 12'h070;
        15'h1F97: data = 12'h070;
        15'h1F98: data = 12'h06E;
        15'h1F99: data = 12'h066;
        15'h1F9A: data = 12'h060;
        15'h1F9B: data = 12'h057;
        15'h1F9C: data = 12'h046;
        15'h1F9D: data = 12'h7BE;
        15'h1F9E: data = 12'h7B0;
        15'h1F9F: data = 12'h7A6;
        15'h1FA0: data = 12'h7A2;
        15'h1FA1: data = 12'h79E;
        15'h1FA2: data = 12'h794;
        15'h1FA3: data = 12'h78F;
        15'h1FA4: data = 12'h77A;
        15'h1FA5: data = 12'h76C;
        15'h1FA6: data = 12'h75B;
        15'h1FA7: data = 12'h746;
        15'h1FA8: data = 12'h734;
        15'h1FA9: data = 12'h72E;
        15'h1FAA: data = 12'h729;
        15'h1FAB: data = 12'h71E;
        15'h1FAC: data = 12'h716;
        15'h1FAD: data = 12'h70F;
        15'h1FAE: data = 12'h6FC;
        15'h1FAF: data = 12'h6E9;
        15'h1FB0: data = 12'h6DE;
        15'h1FB1: data = 12'h6C8;
        15'h1FB2: data = 12'h6B4;
        15'h1FB3: data = 12'h6A4;
        15'h1FB4: data = 12'h696;
        15'h1FB5: data = 12'h688;
        15'h1FB6: data = 12'h682;
        15'h1FB7: data = 12'h673;
        15'h1FB8: data = 12'h668;
        15'h1FB9: data = 12'h65B;
        15'h1FBA: data = 12'h64B;
        15'h1FBB: data = 12'h637;
        15'h1FBC: data = 12'h62A;
        15'h1FBD: data = 12'h60D;
        15'h1FBE: data = 12'h5F8;
        15'h1FBF: data = 12'h5E5;
        15'h1FC0: data = 12'h5CF;
        15'h1FC1: data = 12'h5BE;
        15'h1FC2: data = 12'h5B4;
        15'h1FC3: data = 12'h5A7;
        15'h1FC4: data = 12'h594;
        15'h1FC5: data = 12'h582;
        15'h1FC6: data = 12'h575;
        15'h1FC7: data = 12'h567;
        15'h1FC8: data = 12'h558;
        15'h1FC9: data = 12'h547;
        15'h1FCA: data = 12'h52B;
        15'h1FCB: data = 12'h51D;
        15'h1FCC: data = 12'h507;
        15'h1FCD: data = 12'h4F1;
        15'h1FCE: data = 12'h4D9;
        15'h1FCF: data = 12'h4C7;
        15'h1FD0: data = 12'h4AD;
        15'h1FD1: data = 12'h498;
        15'h1FD2: data = 12'h47F;
        15'h1FD3: data = 12'h469;
        15'h1FD4: data = 12'h450;
        15'h1FD5: data = 12'h442;
        15'h1FD6: data = 12'h42C;
        15'h1FD7: data = 12'h416;
        15'h1FD8: data = 12'h3FE;
        15'h1FD9: data = 12'h3E8;
        15'h1FDA: data = 12'h3D6;
        15'h1FDB: data = 12'h3C1;
        15'h1FDC: data = 12'h3AD;
        15'h1FDD: data = 12'h394;
        15'h1FDE: data = 12'h385;
        15'h1FDF: data = 12'h36C;
        15'h1FE0: data = 12'h35A;
        15'h1FE1: data = 12'h342;
        15'h1FE2: data = 12'h330;
        15'h1FE3: data = 12'h31D;
        15'h1FE4: data = 12'h305;
        15'h1FE5: data = 12'h2EE;
        15'h1FE6: data = 12'h2D8;
        15'h1FE7: data = 12'h2C6;
        15'h1FE8: data = 12'h2AB;
        15'h1FE9: data = 12'h290;
        15'h1FEA: data = 12'h281;
        15'h1FEB: data = 12'h26B;
        15'h1FEC: data = 12'h24F;
        15'h1FED: data = 12'h23A;
        15'h1FEE: data = 12'h21F;
        15'h1FEF: data = 12'h207;
        15'h1FF0: data = 12'h1F7;
        15'h1FF1: data = 12'h1DB;
        15'h1FF2: data = 12'h1C2;
        15'h1FF3: data = 12'h1AC;
        15'h1FF4: data = 12'h194;
        15'h1FF5: data = 12'h17D;
        15'h1FF6: data = 12'h163;
        15'h1FF7: data = 12'h14E;
        15'h1FF8: data = 12'h137;
        15'h1FF9: data = 12'h120;
        15'h1FFA: data = 12'h10D;
        15'h1FFB: data = 12'h0F5;
        15'h1FFC: data = 12'h0DF;
        15'h1FFD: data = 12'h0C5;
        15'h1FFE: data = 12'h0A8;
        15'h1FFF: data = 12'h092;
        15'h2000: data = 12'h07E;
        15'h2001: data = 12'h064;
        15'h2002: data = 12'h04A;
        15'h2003: data = 12'h7E0;
        15'h2004: data = 12'h7D1;
        15'h2005: data = 12'h7BD;
        15'h2006: data = 12'h7A7;
        15'h2007: data = 12'h78F;
        15'h2008: data = 12'h778;
        15'h2009: data = 12'h75D;
        15'h200A: data = 12'h74B;
        15'h200B: data = 12'h735;
        15'h200C: data = 12'h71D;
        15'h200D: data = 12'h708;
        15'h200E: data = 12'h6F0;
        15'h200F: data = 12'h6D8;
        15'h2010: data = 12'h6C3;
        15'h2011: data = 12'h6AC;
        15'h2012: data = 12'h696;
        15'h2013: data = 12'h683;
        15'h2014: data = 12'h668;
        15'h2015: data = 12'h656;
        15'h2016: data = 12'h63C;
        15'h2017: data = 12'h62A;
        15'h2018: data = 12'h610;
        15'h2019: data = 12'h5FA;
        15'h201A: data = 12'h5E1;
        15'h201B: data = 12'h5CD;
        15'h201C: data = 12'h5B9;
        15'h201D: data = 12'h59D;
        15'h201E: data = 12'h58A;
        15'h201F: data = 12'h572;
        15'h2020: data = 12'h55F;
        15'h2021: data = 12'h549;
        15'h2022: data = 12'h533;
        15'h2023: data = 12'h51C;
        15'h2024: data = 12'h508;
        15'h2025: data = 12'h4F3;
        15'h2026: data = 12'h4DC;
        15'h2027: data = 12'h4CB;
        15'h2028: data = 12'h4B8;
        15'h2029: data = 12'h4A7;
        15'h202A: data = 12'h493;
        15'h202B: data = 12'h47F;
        15'h202C: data = 12'h46D;
        15'h202D: data = 12'h459;
        15'h202E: data = 12'h44B;
        15'h202F: data = 12'h43D;
        15'h2030: data = 12'h428;
        15'h2031: data = 12'h41E;
        15'h2032: data = 12'h405;
        15'h2033: data = 12'h3F6;
        15'h2034: data = 12'h3E8;
        15'h2035: data = 12'h3D3;
        15'h2036: data = 12'h3C1;
        15'h2037: data = 12'h3B0;
        15'h2038: data = 12'h39C;
        15'h2039: data = 12'h392;
        15'h203A: data = 12'h376;
        15'h203B: data = 12'h366;
        15'h203C: data = 12'h34F;
        15'h203D: data = 12'h33E;
        15'h203E: data = 12'h330;
        15'h203F: data = 12'h31F;
        15'h2040: data = 12'h30D;
        15'h2041: data = 12'h2FD;
        15'h2042: data = 12'h2F1;
        15'h2043: data = 12'h2E3;
        15'h2044: data = 12'h2D7;
        15'h2045: data = 12'h2D9;
        15'h2046: data = 12'h2C7;
        15'h2047: data = 12'h2BA;
        15'h2048: data = 12'h2AC;
        15'h2049: data = 12'h2A1;
        15'h204A: data = 12'h295;
        15'h204B: data = 12'h283;
        15'h204C: data = 12'h27A;
        15'h204D: data = 12'h268;
        15'h204E: data = 12'h25C;
        15'h204F: data = 12'h248;
        15'h2050: data = 12'h23F;
        15'h2051: data = 12'h22D;
        15'h2052: data = 12'h224;
        15'h2053: data = 12'h217;
        15'h2054: data = 12'h20F;
        15'h2055: data = 12'h20D;
        15'h2056: data = 12'h20A;
        15'h2057: data = 12'h1FA;
        15'h2058: data = 12'h1F9;
        15'h2059: data = 12'h1F2;
        15'h205A: data = 12'h1ED;
        15'h205B: data = 12'h1E3;
        15'h205C: data = 12'h1D5;
        15'h205D: data = 12'h1C8;
        15'h205E: data = 12'h1BF;
        15'h205F: data = 12'h1BB;
        15'h2060: data = 12'h1AF;
        15'h2061: data = 12'h1A3;
        15'h2062: data = 12'h19B;
        15'h2063: data = 12'h194;
        15'h2064: data = 12'h194;
        15'h2065: data = 12'h18F;
        15'h2066: data = 12'h18D;
        15'h2067: data = 12'h189;
        15'h2068: data = 12'h18C;
        15'h2069: data = 12'h186;
        15'h206A: data = 12'h185;
        15'h206B: data = 12'h17C;
        15'h206C: data = 12'h17E;
        15'h206D: data = 12'h172;
        15'h206E: data = 12'h16F;
        15'h206F: data = 12'h16D;
        15'h2070: data = 12'h162;
        15'h2071: data = 12'h15D;
        15'h2072: data = 12'h15C;
        15'h2073: data = 12'h15B;
        15'h2074: data = 12'h158;
        15'h2075: data = 12'h15B;
        15'h2076: data = 12'h15E;
        15'h2077: data = 12'h162;
        15'h2078: data = 12'h164;
        15'h2079: data = 12'h166;
        15'h207A: data = 12'h167;
        15'h207B: data = 12'h16F;
        15'h207C: data = 12'h16F;
        15'h207D: data = 12'h16A;
        15'h207E: data = 12'h167;
        15'h207F: data = 12'h167;
        15'h2080: data = 12'h16A;
        15'h2081: data = 12'h164;
        15'h2082: data = 12'h167;
        15'h2083: data = 12'h16D;
        15'h2084: data = 12'h16E;
        15'h2085: data = 12'h177;
        15'h2086: data = 12'h184;
        15'h2087: data = 12'h187;
        15'h2088: data = 12'h195;
        15'h2089: data = 12'h194;
        15'h208A: data = 12'h19E;
        15'h208B: data = 12'h1A7;
        15'h208C: data = 12'h1AB;
        15'h208D: data = 12'h1B4;
        15'h208E: data = 12'h1AF;
        15'h208F: data = 12'h1B4;
        15'h2090: data = 12'h1B9;
        15'h2091: data = 12'h1BB;
        15'h2092: data = 12'h1BE;
        15'h2093: data = 12'h1C8;
        15'h2094: data = 12'h1D0;
        15'h2095: data = 12'h1DA;
        15'h2096: data = 12'h1E6;
        15'h2097: data = 12'h1F3;
        15'h2098: data = 12'h202;
        15'h2099: data = 12'h20C;
        15'h209A: data = 12'h21D;
        15'h209B: data = 12'h220;
        15'h209C: data = 12'h231;
        15'h209D: data = 12'h239;
        15'h209E: data = 12'h246;
        15'h209F: data = 12'h24D;
        15'h20A0: data = 12'h25A;
        15'h20A1: data = 12'h25C;
        15'h20A2: data = 12'h26A;
        15'h20A3: data = 12'h26B;
        15'h20A4: data = 12'h27B;
        15'h20A5: data = 12'h287;
        15'h20A6: data = 12'h290;
        15'h20A7: data = 12'h2A1;
        15'h20A8: data = 12'h2B1;
        15'h20A9: data = 12'h2C2;
        15'h20AA: data = 12'h2D1;
        15'h20AB: data = 12'h2DE;
        15'h20AC: data = 12'h2F3;
        15'h20AD: data = 12'h305;
        15'h20AE: data = 12'h317;
        15'h20AF: data = 12'h328;
        15'h20B0: data = 12'h337;
        15'h20B1: data = 12'h344;
        15'h20B2: data = 12'h354;
        15'h20B3: data = 12'h364;
        15'h20B4: data = 12'h370;
        15'h20B5: data = 12'h37B;
        15'h20B6: data = 12'h38F;
        15'h20B7: data = 12'h395;
        15'h20B8: data = 12'h3A8;
        15'h20B9: data = 12'h3B5;
        15'h20BA: data = 12'h3C5;
        15'h20BB: data = 12'h3DD;
        15'h20BC: data = 12'h3EF;
        15'h20BD: data = 12'h3FD;
        15'h20BE: data = 12'h418;
        15'h20BF: data = 12'h42D;
        15'h20C0: data = 12'h443;
        15'h20C1: data = 12'h459;
        15'h20C2: data = 12'h46C;
        15'h20C3: data = 12'h481;
        15'h20C4: data = 12'h493;
        15'h20C5: data = 12'h4AC;
        15'h20C6: data = 12'h4BA;
        15'h20C7: data = 12'h4D1;
        15'h20C8: data = 12'h4E3;
        15'h20C9: data = 12'h4F4;
        15'h20CA: data = 12'h507;
        15'h20CB: data = 12'h516;
        15'h20CC: data = 12'h525;
        15'h20CD: data = 12'h53C;
        15'h20CE: data = 12'h550;
        15'h20CF: data = 12'h562;
        15'h20D0: data = 12'h573;
        15'h20D1: data = 12'h58B;
        15'h20D2: data = 12'h5A0;
        15'h20D3: data = 12'h5BC;
        15'h20D4: data = 12'h5CD;
        15'h20D5: data = 12'h5E7;
        15'h20D6: data = 12'h605;
        15'h20D7: data = 12'h61C;
        15'h20D8: data = 12'h632;
        15'h20D9: data = 12'h64B;
        15'h20DA: data = 12'h661;
        15'h20DB: data = 12'h676;
        15'h20DC: data = 12'h693;
        15'h20DD: data = 12'h6A1;
        15'h20DE: data = 12'h6B8;
        15'h20DF: data = 12'h6CB;
        15'h20E0: data = 12'h6E1;
        15'h20E1: data = 12'h6F6;
        15'h20E2: data = 12'h70A;
        15'h20E3: data = 12'h71F;
        15'h20E4: data = 12'h735;
        15'h20E5: data = 12'h743;
        15'h20E6: data = 12'h75C;
        15'h20E7: data = 12'h771;
        15'h20E8: data = 12'h78D;
        15'h20E9: data = 12'h7A1;
        15'h20EA: data = 12'h7B8;
        15'h20EB: data = 12'h7D6;
        15'h20EC: data = 12'h7E9;
        15'h20ED: data = 12'h804;
        15'h20EE: data = 12'h073;
        15'h20EF: data = 12'h08C;
        15'h20F0: data = 12'h0A1;
        15'h20F1: data = 12'h0B4;
        15'h20F2: data = 12'h0D2;
        15'h20F3: data = 12'h0EC;
        15'h20F4: data = 12'h0FE;
        15'h20F5: data = 12'h115;
        15'h20F6: data = 12'h12B;
        15'h20F7: data = 12'h141;
        15'h20F8: data = 12'h154;
        15'h20F9: data = 12'h16C;
        15'h20FA: data = 12'h17E;
        15'h20FB: data = 12'h197;
        15'h20FC: data = 12'h1B0;
        15'h20FD: data = 12'h1BC;
        15'h20FE: data = 12'h1D7;
        15'h20FF: data = 12'h1EC;
        15'h2100: data = 12'h202;
        15'h2101: data = 12'h216;
        15'h2102: data = 12'h22E;
        15'h2103: data = 12'h24A;
        15'h2104: data = 12'h25F;
        15'h2105: data = 12'h277;
        15'h2106: data = 12'h28C;
        15'h2107: data = 12'h2A6;
        15'h2108: data = 12'h2BD;
        15'h2109: data = 12'h2D2;
        15'h210A: data = 12'h2F1;
        15'h210B: data = 12'h306;
        15'h210C: data = 12'h321;
        15'h210D: data = 12'h337;
        15'h210E: data = 12'h34D;
        15'h210F: data = 12'h368;
        15'h2110: data = 12'h37D;
        15'h2111: data = 12'h398;
        15'h2112: data = 12'h3AB;
        15'h2113: data = 12'h3C3;
        15'h2114: data = 12'h3DD;
        15'h2115: data = 12'h3F2;
        15'h2116: data = 12'h400;
        15'h2117: data = 12'h418;
        15'h2118: data = 12'h42D;
        15'h2119: data = 12'h442;
        15'h211A: data = 12'h450;
        15'h211B: data = 12'h464;
        15'h211C: data = 12'h47E;
        15'h211D: data = 12'h493;
        15'h211E: data = 12'h4A7;
        15'h211F: data = 12'h4B7;
        15'h2120: data = 12'h4C6;
        15'h2121: data = 12'h4DA;
        15'h2122: data = 12'h4EE;
        15'h2123: data = 12'h507;
        15'h2124: data = 12'h511;
        15'h2125: data = 12'h523;
        15'h2126: data = 12'h53A;
        15'h2127: data = 12'h548;
        15'h2128: data = 12'h55B;
        15'h2129: data = 12'h569;
        15'h212A: data = 12'h57E;
        15'h212B: data = 12'h590;
        15'h212C: data = 12'h5A5;
        15'h212D: data = 12'h5B9;
        15'h212E: data = 12'h5C8;
        15'h212F: data = 12'h5D8;
        15'h2130: data = 12'h5EB;
        15'h2131: data = 12'h5FE;
        15'h2132: data = 12'h60C;
        15'h2133: data = 12'h61B;
        15'h2134: data = 12'h62D;
        15'h2135: data = 12'h63B;
        15'h2136: data = 12'h64F;
        15'h2137: data = 12'h663;
        15'h2138: data = 12'h675;
        15'h2139: data = 12'h685;
        15'h213A: data = 12'h698;
        15'h213B: data = 12'h6A4;
        15'h213C: data = 12'h6B5;
        15'h213D: data = 12'h6C6;
        15'h213E: data = 12'h6D3;
        15'h213F: data = 12'h6DD;
        15'h2140: data = 12'h6EF;
        15'h2141: data = 12'h700;
        15'h2142: data = 12'h708;
        15'h2143: data = 12'h716;
        15'h2144: data = 12'h723;
        15'h2145: data = 12'h734;
        15'h2146: data = 12'h73A;
        15'h2147: data = 12'h743;
        15'h2148: data = 12'h750;
        15'h2149: data = 12'h75E;
        15'h214A: data = 12'h769;
        15'h214B: data = 12'h775;
        15'h214C: data = 12'h77D;
        15'h214D: data = 12'h78A;
        15'h214E: data = 12'h791;
        15'h214F: data = 12'h79B;
        15'h2150: data = 12'h7A2;
        15'h2151: data = 12'h7AC;
        15'h2152: data = 12'h7B7;
        15'h2153: data = 12'h7BC;
        15'h2154: data = 12'h7C6;
        15'h2155: data = 12'h7CD;
        15'h2156: data = 12'h7D6;
        15'h2157: data = 12'h7DC;
        15'h2158: data = 12'h7E6;
        15'h2159: data = 12'h7E9;
        15'h215A: data = 12'h7ED;
        15'h215B: data = 12'h7F7;
        15'h215C: data = 12'h7FE;
        15'h215D: data = 12'h7FF;
        15'h215E: data = 12'h802;
        15'h215F: data = 12'h80B;
        15'h2160: data = 12'h766;
        15'h2161: data = 12'h086;
        15'h2162: data = 12'h094;
        15'h2163: data = 12'h097;
        15'h2164: data = 12'h098;
        15'h2165: data = 12'h09D;
        15'h2166: data = 12'h0A3;
        15'h2167: data = 12'h0AB;
        15'h2168: data = 12'h0AD;
        15'h2169: data = 12'h0AC;
        15'h216A: data = 12'h0B6;
        15'h216B: data = 12'h0BB;
        15'h216C: data = 12'h0B9;
        15'h216D: data = 12'h0BA;
        15'h216E: data = 12'h0C8;
        15'h216F: data = 12'h0C9;
        15'h2170: data = 12'h0CE;
        15'h2171: data = 12'h0D0;
        15'h2172: data = 12'h0D3;
        15'h2173: data = 12'h0D2;
        15'h2174: data = 12'h0D6;
        15'h2175: data = 12'h0CD;
        15'h2176: data = 12'h0D0;
        15'h2177: data = 12'h0CD;
        15'h2178: data = 12'h0CB;
        15'h2179: data = 12'h0C8;
        15'h217A: data = 12'h0BF;
        15'h217B: data = 12'h0B6;
        15'h217C: data = 12'h0AD;
        15'h217D: data = 12'h0AD;
        15'h217E: data = 12'h0A6;
        15'h217F: data = 12'h0A8;
        15'h2180: data = 12'h0A9;
        15'h2181: data = 12'h0AF;
        15'h2182: data = 12'h0AD;
        15'h2183: data = 12'h0A2;
        15'h2184: data = 12'h0A7;
        15'h2185: data = 12'h09D;
        15'h2186: data = 12'h092;
        15'h2187: data = 12'h083;
        15'h2188: data = 12'h075;
        15'h2189: data = 12'h074;
        15'h218A: data = 12'h06B;
        15'h218B: data = 12'h069;
        15'h218C: data = 12'h067;
        15'h218D: data = 12'h066;
        15'h218E: data = 12'h05D;
        15'h218F: data = 12'h057;
        15'h2190: data = 12'h04C;
        15'h2191: data = 12'h038;
        15'h2192: data = 12'h7B9;
        15'h2193: data = 12'h7A9;
        15'h2194: data = 12'h7A2;
        15'h2195: data = 12'h797;
        15'h2196: data = 12'h791;
        15'h2197: data = 12'h78F;
        15'h2198: data = 12'h780;
        15'h2199: data = 12'h774;
        15'h219A: data = 12'h760;
        15'h219B: data = 12'h74C;
        15'h219C: data = 12'h73A;
        15'h219D: data = 12'h72E;
        15'h219E: data = 12'h723;
        15'h219F: data = 12'h71B;
        15'h21A0: data = 12'h714;
        15'h21A1: data = 12'h70B;
        15'h21A2: data = 12'h6FF;
        15'h21A3: data = 12'h6EA;
        15'h21A4: data = 12'h6E1;
        15'h21A5: data = 12'h6CA;
        15'h21A6: data = 12'h6B8;
        15'h21A7: data = 12'h6A7;
        15'h21A8: data = 12'h697;
        15'h21A9: data = 12'h686;
        15'h21AA: data = 12'h67D;
        15'h21AB: data = 12'h674;
        15'h21AC: data = 12'h669;
        15'h21AD: data = 12'h65B;
        15'h21AE: data = 12'h647;
        15'h21AF: data = 12'h638;
        15'h21B0: data = 12'h62E;
        15'h21B1: data = 12'h610;
        15'h21B2: data = 12'h5FA;
        15'h21B3: data = 12'h5EA;
        15'h21B4: data = 12'h5CF;
        15'h21B5: data = 12'h5BF;
        15'h21B6: data = 12'h5B1;
        15'h21B7: data = 12'h5A4;
        15'h21B8: data = 12'h58F;
        15'h21B9: data = 12'h581;
        15'h21BA: data = 12'h56F;
        15'h21BB: data = 12'h563;
        15'h21BC: data = 12'h554;
        15'h21BD: data = 12'h544;
        15'h21BE: data = 12'h52E;
        15'h21BF: data = 12'h51D;
        15'h21C0: data = 12'h509;
        15'h21C1: data = 12'h4F3;
        15'h21C2: data = 12'h4DA;
        15'h21C3: data = 12'h4C5;
        15'h21C4: data = 12'h4AF;
        15'h21C5: data = 12'h49A;
        15'h21C6: data = 12'h481;
        15'h21C7: data = 12'h469;
        15'h21C8: data = 12'h451;
        15'h21C9: data = 12'h441;
        15'h21CA: data = 12'h42C;
        15'h21CB: data = 12'h416;
        15'h21CC: data = 12'h3FF;
        15'h21CD: data = 12'h3E7;
        15'h21CE: data = 12'h3D5;
        15'h21CF: data = 12'h3C4;
        15'h21D0: data = 12'h3B1;
        15'h21D1: data = 12'h395;
        15'h21D2: data = 12'h384;
        15'h21D3: data = 12'h36C;
        15'h21D4: data = 12'h35B;
        15'h21D5: data = 12'h346;
        15'h21D6: data = 12'h32F;
        15'h21D7: data = 12'h31F;
        15'h21D8: data = 12'h302;
        15'h21D9: data = 12'h2F2;
        15'h21DA: data = 12'h2DD;
        15'h21DB: data = 12'h2C7;
        15'h21DC: data = 12'h2AB;
        15'h21DD: data = 12'h292;
        15'h21DE: data = 12'h281;
        15'h21DF: data = 12'h26B;
        15'h21E0: data = 12'h24F;
        15'h21E1: data = 12'h23B;
        15'h21E2: data = 12'h21F;
        15'h21E3: data = 12'h20C;
        15'h21E4: data = 12'h1F5;
        15'h21E5: data = 12'h1DA;
        15'h21E6: data = 12'h1C1;
        15'h21E7: data = 12'h1AA;
        15'h21E8: data = 12'h193;
        15'h21E9: data = 12'h17F;
        15'h21EA: data = 12'h167;
        15'h21EB: data = 12'h14F;
        15'h21EC: data = 12'h13B;
        15'h21ED: data = 12'h121;
        15'h21EE: data = 12'h107;
        15'h21EF: data = 12'h0F2;
        15'h21F0: data = 12'h0DF;
        15'h21F1: data = 12'h0C1;
        15'h21F2: data = 12'h0A6;
        15'h21F3: data = 12'h08F;
        15'h21F4: data = 12'h081;
        15'h21F5: data = 12'h065;
        15'h21F6: data = 12'h04D;
        15'h21F7: data = 12'h7E2;
        15'h21F8: data = 12'h7CF;
        15'h21F9: data = 12'h7BC;
        15'h21FA: data = 12'h7A6;
        15'h21FB: data = 12'h78D;
        15'h21FC: data = 12'h773;
        15'h21FD: data = 12'h75E;
        15'h21FE: data = 12'h74A;
        15'h21FF: data = 12'h734;
        15'h2200: data = 12'h71E;
        15'h2201: data = 12'h709;
        15'h2202: data = 12'h6ED;
        15'h2203: data = 12'h6D6;
        15'h2204: data = 12'h6C3;
        15'h2205: data = 12'h6AD;
        15'h2206: data = 12'h696;
        15'h2207: data = 12'h686;
        15'h2208: data = 12'h667;
        15'h2209: data = 12'h655;
        15'h220A: data = 12'h63B;
        15'h220B: data = 12'h62A;
        15'h220C: data = 12'h614;
        15'h220D: data = 12'h5F9;
        15'h220E: data = 12'h5E1;
        15'h220F: data = 12'h5CC;
        15'h2210: data = 12'h5BB;
        15'h2211: data = 12'h59D;
        15'h2212: data = 12'h585;
        15'h2213: data = 12'h571;
        15'h2214: data = 12'h55F;
        15'h2215: data = 12'h547;
        15'h2216: data = 12'h533;
        15'h2217: data = 12'h51A;
        15'h2218: data = 12'h50A;
        15'h2219: data = 12'h4F3;
        15'h221A: data = 12'h4DC;
        15'h221B: data = 12'h4CB;
        15'h221C: data = 12'h4B5;
        15'h221D: data = 12'h4A4;
        15'h221E: data = 12'h492;
        15'h221F: data = 12'h47C;
        15'h2220: data = 12'h46E;
        15'h2221: data = 12'h457;
        15'h2222: data = 12'h44B;
        15'h2223: data = 12'h43D;
        15'h2224: data = 12'h42A;
        15'h2225: data = 12'h418;
        15'h2226: data = 12'h408;
        15'h2227: data = 12'h3F8;
        15'h2228: data = 12'h3EB;
        15'h2229: data = 12'h3D4;
        15'h222A: data = 12'h3BE;
        15'h222B: data = 12'h3B0;
        15'h222C: data = 12'h39C;
        15'h222D: data = 12'h391;
        15'h222E: data = 12'h377;
        15'h222F: data = 12'h365;
        15'h2230: data = 12'h353;
        15'h2231: data = 12'h341;
        15'h2232: data = 12'h32E;
        15'h2233: data = 12'h31F;
        15'h2234: data = 12'h30E;
        15'h2235: data = 12'h2FF;
        15'h2236: data = 12'h2F1;
        15'h2237: data = 12'h2E3;
        15'h2238: data = 12'h2D4;
        15'h2239: data = 12'h2D3;
        15'h223A: data = 12'h2C9;
        15'h223B: data = 12'h2BB;
        15'h223C: data = 12'h2AF;
        15'h223D: data = 12'h2A3;
        15'h223E: data = 12'h294;
        15'h223F: data = 12'h284;
        15'h2240: data = 12'h27B;
        15'h2241: data = 12'h269;
        15'h2242: data = 12'h260;
        15'h2243: data = 12'h24A;
        15'h2244: data = 12'h241;
        15'h2245: data = 12'h230;
        15'h2246: data = 12'h226;
        15'h2247: data = 12'h218;
        15'h2248: data = 12'h212;
        15'h2249: data = 12'h209;
        15'h224A: data = 12'h206;
        15'h224B: data = 12'h1FE;
        15'h224C: data = 12'h1F8;
        15'h224D: data = 12'h1F4;
        15'h224E: data = 12'h1EB;
        15'h224F: data = 12'h1E1;
        15'h2250: data = 12'h1D7;
        15'h2251: data = 12'h1CB;
        15'h2252: data = 12'h1C2;
        15'h2253: data = 12'h1BF;
        15'h2254: data = 12'h1AF;
        15'h2255: data = 12'h1A9;
        15'h2256: data = 12'h19D;
        15'h2257: data = 12'h194;
        15'h2258: data = 12'h193;
        15'h2259: data = 12'h18F;
        15'h225A: data = 12'h18A;
        15'h225B: data = 12'h18E;
        15'h225C: data = 12'h18D;
        15'h225D: data = 12'h188;
        15'h225E: data = 12'h189;
        15'h225F: data = 12'h180;
        15'h2260: data = 12'h182;
        15'h2261: data = 12'h176;
        15'h2262: data = 12'h173;
        15'h2263: data = 12'h170;
        15'h2264: data = 12'h164;
        15'h2265: data = 12'h15F;
        15'h2266: data = 12'h15E;
        15'h2267: data = 12'h15D;
        15'h2268: data = 12'h159;
        15'h2269: data = 12'h159;
        15'h226A: data = 12'h15F;
        15'h226B: data = 12'h163;
        15'h226C: data = 12'h164;
        15'h226D: data = 12'h168;
        15'h226E: data = 12'h169;
        15'h226F: data = 12'h172;
        15'h2270: data = 12'h16E;
        15'h2271: data = 12'h16C;
        15'h2272: data = 12'h16B;
        15'h2273: data = 12'h167;
        15'h2274: data = 12'h16B;
        15'h2275: data = 12'h168;
        15'h2276: data = 12'h16A;
        15'h2277: data = 12'h16E;
        15'h2278: data = 12'h16E;
        15'h2279: data = 12'h178;
        15'h227A: data = 12'h184;
        15'h227B: data = 12'h184;
        15'h227C: data = 12'h192;
        15'h227D: data = 12'h192;
        15'h227E: data = 12'h19E;
        15'h227F: data = 12'h1A5;
        15'h2280: data = 12'h1AB;
        15'h2281: data = 12'h1B1;
        15'h2282: data = 12'h1B4;
        15'h2283: data = 12'h1B7;
        15'h2284: data = 12'h1B9;
        15'h2285: data = 12'h1C0;
        15'h2286: data = 12'h1C4;
        15'h2287: data = 12'h1CB;
        15'h2288: data = 12'h1D0;
        15'h2289: data = 12'h1DC;
        15'h228A: data = 12'h1E4;
        15'h228B: data = 12'h1F5;
        15'h228C: data = 12'h1FE;
        15'h228D: data = 12'h20B;
        15'h228E: data = 12'h21E;
        15'h228F: data = 12'h224;
        15'h2290: data = 12'h234;
        15'h2291: data = 12'h23C;
        15'h2292: data = 12'h245;
        15'h2293: data = 12'h24D;
        15'h2294: data = 12'h25A;
        15'h2295: data = 12'h25F;
        15'h2296: data = 12'h268;
        15'h2297: data = 12'h26E;
        15'h2298: data = 12'h27D;
        15'h2299: data = 12'h287;
        15'h229A: data = 12'h291;
        15'h229B: data = 12'h29E;
        15'h229C: data = 12'h2B2;
        15'h229D: data = 12'h2C1;
        15'h229E: data = 12'h2D2;
        15'h229F: data = 12'h2DE;
        15'h22A0: data = 12'h2F4;
        15'h22A1: data = 12'h304;
        15'h22A2: data = 12'h318;
        15'h22A3: data = 12'h329;
        15'h22A4: data = 12'h335;
        15'h22A5: data = 12'h346;
        15'h22A6: data = 12'h351;
        15'h22A7: data = 12'h362;
        15'h22A8: data = 12'h370;
        15'h22A9: data = 12'h37E;
        15'h22AA: data = 12'h391;
        15'h22AB: data = 12'h394;
        15'h22AC: data = 12'h3AA;
        15'h22AD: data = 12'h3BB;
        15'h22AE: data = 12'h3C4;
        15'h22AF: data = 12'h3DD;
        15'h22B0: data = 12'h3EB;
        15'h22B1: data = 12'h3FC;
        15'h22B2: data = 12'h415;
        15'h22B3: data = 12'h42C;
        15'h22B4: data = 12'h444;
        15'h22B5: data = 12'h457;
        15'h22B6: data = 12'h46B;
        15'h22B7: data = 12'h481;
        15'h22B8: data = 12'h493;
        15'h22B9: data = 12'h4A9;
        15'h22BA: data = 12'h4B8;
        15'h22BB: data = 12'h4CF;
        15'h22BC: data = 12'h4E1;
        15'h22BD: data = 12'h4F3;
        15'h22BE: data = 12'h509;
        15'h22BF: data = 12'h517;
        15'h22C0: data = 12'h525;
        15'h22C1: data = 12'h539;
        15'h22C2: data = 12'h54F;
        15'h22C3: data = 12'h562;
        15'h22C4: data = 12'h574;
        15'h22C5: data = 12'h58B;
        15'h22C6: data = 12'h5A2;
        15'h22C7: data = 12'h5B9;
        15'h22C8: data = 12'h5CF;
        15'h22C9: data = 12'h5E3;
        15'h22CA: data = 12'h601;
        15'h22CB: data = 12'h61B;
        15'h22CC: data = 12'h630;
        15'h22CD: data = 12'h646;
        15'h22CE: data = 12'h662;
        15'h22CF: data = 12'h677;
        15'h22D0: data = 12'h692;
        15'h22D1: data = 12'h6A0;
        15'h22D2: data = 12'h6B5;
        15'h22D3: data = 12'h6D1;
        15'h22D4: data = 12'h6E1;
        15'h22D5: data = 12'h6F8;
        15'h22D6: data = 12'h70B;
        15'h22D7: data = 12'h71F;
        15'h22D8: data = 12'h738;
        15'h22D9: data = 12'h745;
        15'h22DA: data = 12'h75C;
        15'h22DB: data = 12'h773;
        15'h22DC: data = 12'h78E;
        15'h22DD: data = 12'h79F;
        15'h22DE: data = 12'h7BB;
        15'h22DF: data = 12'h7D6;
        15'h22E0: data = 12'h7EC;
        15'h22E1: data = 12'h806;
        15'h22E2: data = 12'h073;
        15'h22E3: data = 12'h08E;
        15'h22E4: data = 12'h0A1;
        15'h22E5: data = 12'h0B7;
        15'h22E6: data = 12'h0D1;
        15'h22E7: data = 12'h0EA;
        15'h22E8: data = 12'h100;
        15'h22E9: data = 12'h115;
        15'h22EA: data = 12'h129;
        15'h22EB: data = 12'h140;
        15'h22EC: data = 12'h157;
        15'h22ED: data = 12'h16C;
        15'h22EE: data = 12'h183;
        15'h22EF: data = 12'h198;
        15'h22F0: data = 12'h1B2;
        15'h22F1: data = 12'h1C0;
        15'h22F2: data = 12'h1D8;
        15'h22F3: data = 12'h1F0;
        15'h22F4: data = 12'h208;
        15'h22F5: data = 12'h215;
        15'h22F6: data = 12'h234;
        15'h22F7: data = 12'h249;
        15'h22F8: data = 12'h261;
        15'h22F9: data = 12'h276;
        15'h22FA: data = 12'h289;
        15'h22FB: data = 12'h2A7;
        15'h22FC: data = 12'h2C2;
        15'h22FD: data = 12'h2D4;
        15'h22FE: data = 12'h2F0;
        15'h22FF: data = 12'h30B;
        15'h2300: data = 12'h323;
        15'h2301: data = 12'h336;
        15'h2302: data = 12'h34E;
        15'h2303: data = 12'h369;
        15'h2304: data = 12'h37D;
        15'h2305: data = 12'h39B;
        15'h2306: data = 12'h3AB;
        15'h2307: data = 12'h3C2;
        15'h2308: data = 12'h3DC;
        15'h2309: data = 12'h3F2;
        15'h230A: data = 12'h403;
        15'h230B: data = 12'h417;
        15'h230C: data = 12'h430;
        15'h230D: data = 12'h447;
        15'h230E: data = 12'h454;
        15'h230F: data = 12'h467;
        15'h2310: data = 12'h47F;
        15'h2311: data = 12'h496;
        15'h2312: data = 12'h4A9;
        15'h2313: data = 12'h4B9;
        15'h2314: data = 12'h4C9;
        15'h2315: data = 12'h4DE;
        15'h2316: data = 12'h4F2;
        15'h2317: data = 12'h507;
        15'h2318: data = 12'h512;
        15'h2319: data = 12'h525;
        15'h231A: data = 12'h53E;
        15'h231B: data = 12'h549;
        15'h231C: data = 12'h55D;
        15'h231D: data = 12'h56B;
        15'h231E: data = 12'h581;
        15'h231F: data = 12'h593;
        15'h2320: data = 12'h5A5;
        15'h2321: data = 12'h5B9;
        15'h2322: data = 12'h5C4;
        15'h2323: data = 12'h5D7;
        15'h2324: data = 12'h5ED;
        15'h2325: data = 12'h5FD;
        15'h2326: data = 12'h60F;
        15'h2327: data = 12'h61E;
        15'h2328: data = 12'h62C;
        15'h2329: data = 12'h63C;
        15'h232A: data = 12'h651;
        15'h232B: data = 12'h663;
        15'h232C: data = 12'h672;
        15'h232D: data = 12'h682;
        15'h232E: data = 12'h695;
        15'h232F: data = 12'h6A5;
        15'h2330: data = 12'h6B2;
        15'h2331: data = 12'h6C6;
        15'h2332: data = 12'h6D2;
        15'h2333: data = 12'h6DC;
        15'h2334: data = 12'h6EC;
        15'h2335: data = 12'h6F9;
        15'h2336: data = 12'h70A;
        15'h2337: data = 12'h715;
        15'h2338: data = 12'h727;
        15'h2339: data = 12'h734;
        15'h233A: data = 12'h737;
        15'h233B: data = 12'h745;
        15'h233C: data = 12'h74F;
        15'h233D: data = 12'h760;
        15'h233E: data = 12'h766;
        15'h233F: data = 12'h777;
        15'h2340: data = 12'h77F;
        15'h2341: data = 12'h78C;
        15'h2342: data = 12'h796;
        15'h2343: data = 12'h79E;
        15'h2344: data = 12'h7A5;
        15'h2345: data = 12'h7B0;
        15'h2346: data = 12'h7B8;
        15'h2347: data = 12'h7C0;
        15'h2348: data = 12'h7C5;
        15'h2349: data = 12'h7CC;
        15'h234A: data = 12'h7D4;
        15'h234B: data = 12'h7DC;
        15'h234C: data = 12'h7E8;
        15'h234D: data = 12'h7EB;
        15'h234E: data = 12'h7F2;
        15'h234F: data = 12'h7F9;
        15'h2350: data = 12'h7FE;
        15'h2351: data = 12'h802;
        15'h2352: data = 12'h804;
        15'h2353: data = 12'h80B;
        15'h2354: data = 12'h790;
        15'h2355: data = 12'h089;
        15'h2356: data = 12'h093;
        15'h2357: data = 12'h097;
        15'h2358: data = 12'h09E;
        15'h2359: data = 12'h0A2;
        15'h235A: data = 12'h0A2;
        15'h235B: data = 12'h0A9;
        15'h235C: data = 12'h0AA;
        15'h235D: data = 12'h0AC;
        15'h235E: data = 12'h0B8;
        15'h235F: data = 12'h0B7;
        15'h2360: data = 12'h0B9;
        15'h2361: data = 12'h0BC;
        15'h2362: data = 12'h0C7;
        15'h2363: data = 12'h0C8;
        15'h2364: data = 12'h0C9;
        15'h2365: data = 12'h0CD;
        15'h2366: data = 12'h0D1;
        15'h2367: data = 12'h0D5;
        15'h2368: data = 12'h0D6;
        15'h2369: data = 12'h0CE;
        15'h236A: data = 12'h0CB;
        15'h236B: data = 12'h0CE;
        15'h236C: data = 12'h0CB;
        15'h236D: data = 12'h0CA;
        15'h236E: data = 12'h0BE;
        15'h236F: data = 12'h0BA;
        15'h2370: data = 12'h0AD;
        15'h2371: data = 12'h0B1;
        15'h2372: data = 12'h0A8;
        15'h2373: data = 12'h0AA;
        15'h2374: data = 12'h0AA;
        15'h2375: data = 12'h0AE;
        15'h2376: data = 12'h0AF;
        15'h2377: data = 12'h0A8;
        15'h2378: data = 12'h0A7;
        15'h2379: data = 12'h09D;
        15'h237A: data = 12'h090;
        15'h237B: data = 12'h083;
        15'h237C: data = 12'h075;
        15'h237D: data = 12'h072;
        15'h237E: data = 12'h06D;
        15'h237F: data = 12'h068;
        15'h2380: data = 12'h066;
        15'h2381: data = 12'h066;
        15'h2382: data = 12'h05F;
        15'h2383: data = 12'h059;
        15'h2384: data = 12'h04B;
        15'h2385: data = 12'h03A;
        15'h2386: data = 12'h7BA;
        15'h2387: data = 12'h7A8;
        15'h2388: data = 12'h7A2;
        15'h2389: data = 12'h79A;
        15'h238A: data = 12'h791;
        15'h238B: data = 12'h78E;
        15'h238C: data = 12'h780;
        15'h238D: data = 12'h771;
        15'h238E: data = 12'h760;
        15'h238F: data = 12'h74B;
        15'h2390: data = 12'h738;
        15'h2391: data = 12'h730;
        15'h2392: data = 12'h724;
        15'h2393: data = 12'h71B;
        15'h2394: data = 12'h714;
        15'h2395: data = 12'h70A;
        15'h2396: data = 12'h6FD;
        15'h2397: data = 12'h6EB;
        15'h2398: data = 12'h6DD;
        15'h2399: data = 12'h6CA;
        15'h239A: data = 12'h6B6;
        15'h239B: data = 12'h6A9;
        15'h239C: data = 12'h696;
        15'h239D: data = 12'h687;
        15'h239E: data = 12'h67A;
        15'h239F: data = 12'h672;
        15'h23A0: data = 12'h666;
        15'h23A1: data = 12'h65B;
        15'h23A2: data = 12'h648;
        15'h23A3: data = 12'h636;
        15'h23A4: data = 12'h62B;
        15'h23A5: data = 12'h60D;
        15'h23A6: data = 12'h5FA;
        15'h23A7: data = 12'h5E9;
        15'h23A8: data = 12'h5D1;
        15'h23A9: data = 12'h5C0;
        15'h23AA: data = 12'h5B2;
        15'h23AB: data = 12'h5A4;
        15'h23AC: data = 12'h590;
        15'h23AD: data = 12'h585;
        15'h23AE: data = 12'h56E;
        15'h23AF: data = 12'h565;
        15'h23B0: data = 12'h557;
        15'h23B1: data = 12'h544;
        15'h23B2: data = 12'h52E;
        15'h23B3: data = 12'h51D;
        15'h23B4: data = 12'h507;
        15'h23B5: data = 12'h4F5;
        15'h23B6: data = 12'h4D9;
        15'h23B7: data = 12'h4C5;
        15'h23B8: data = 12'h4B0;
        15'h23B9: data = 12'h496;
        15'h23BA: data = 12'h483;
        15'h23BB: data = 12'h469;
        15'h23BC: data = 12'h44F;
        15'h23BD: data = 12'h440;
        15'h23BE: data = 12'h42A;
        15'h23BF: data = 12'h414;
        15'h23C0: data = 12'h403;
        15'h23C1: data = 12'h3E7;
        15'h23C2: data = 12'h3D6;
        15'h23C3: data = 12'h3C3;
        15'h23C4: data = 12'h3B0;
        15'h23C5: data = 12'h397;
        15'h23C6: data = 12'h384;
        15'h23C7: data = 12'h36E;
        15'h23C8: data = 12'h357;
        15'h23C9: data = 12'h343;
        15'h23CA: data = 12'h334;
        15'h23CB: data = 12'h31B;
        15'h23CC: data = 12'h302;
        15'h23CD: data = 12'h2F0;
        15'h23CE: data = 12'h2DF;
        15'h23CF: data = 12'h2C5;
        15'h23D0: data = 12'h2AD;
        15'h23D1: data = 12'h291;
        15'h23D2: data = 12'h282;
        15'h23D3: data = 12'h269;
        15'h23D4: data = 12'h250;
        15'h23D5: data = 12'h239;
        15'h23D6: data = 12'h21E;
        15'h23D7: data = 12'h20C;
        15'h23D8: data = 12'h1F9;
        15'h23D9: data = 12'h1DC;
        15'h23DA: data = 12'h1C1;
        15'h23DB: data = 12'h1AB;
        15'h23DC: data = 12'h196;
        15'h23DD: data = 12'h180;
        15'h23DE: data = 12'h167;
        15'h23DF: data = 12'h150;
        15'h23E0: data = 12'h139;
        15'h23E1: data = 12'h121;
        15'h23E2: data = 12'h109;
        15'h23E3: data = 12'h0F3;
        15'h23E4: data = 12'h0DB;
        15'h23E5: data = 12'h0C2;
        15'h23E6: data = 12'h0AB;
        15'h23E7: data = 12'h093;
        15'h23E8: data = 12'h07F;
        15'h23E9: data = 12'h063;
        15'h23EA: data = 12'h050;
        15'h23EB: data = 12'h7DF;
        15'h23EC: data = 12'h7D0;
        15'h23ED: data = 12'h7BD;
        15'h23EE: data = 12'h7A1;
        15'h23EF: data = 12'h78B;
        15'h23F0: data = 12'h777;
        15'h23F1: data = 12'h75E;
        15'h23F2: data = 12'h74B;
        15'h23F3: data = 12'h734;
        15'h23F4: data = 12'h71C;
        15'h23F5: data = 12'h709;
        15'h23F6: data = 12'h6F0;
        15'h23F7: data = 12'h6DB;
        15'h23F8: data = 12'h6C5;
        15'h23F9: data = 12'h6AC;
        15'h23FA: data = 12'h696;
        15'h23FB: data = 12'h683;
        15'h23FC: data = 12'h668;
        15'h23FD: data = 12'h655;
        15'h23FE: data = 12'h63D;
        15'h23FF: data = 12'h62C;
        15'h2400: data = 12'h616;
        15'h2401: data = 12'h5F9;
        15'h2402: data = 12'h5E4;
        15'h2403: data = 12'h5CB;
        15'h2404: data = 12'h5BA;
        15'h2405: data = 12'h59D;
        15'h2406: data = 12'h588;
        15'h2407: data = 12'h572;
        15'h2408: data = 12'h55E;
        15'h2409: data = 12'h548;
        15'h240A: data = 12'h530;
        15'h240B: data = 12'h518;
        15'h240C: data = 12'h509;
        15'h240D: data = 12'h4EF;
        15'h240E: data = 12'h4DC;
        15'h240F: data = 12'h4C9;
        15'h2410: data = 12'h4B7;
        15'h2411: data = 12'h4A6;
        15'h2412: data = 12'h491;
        15'h2413: data = 12'h47F;
        15'h2414: data = 12'h46D;
        15'h2415: data = 12'h45A;
        15'h2416: data = 12'h44B;
        15'h2417: data = 12'h43E;
        15'h2418: data = 12'h429;
        15'h2419: data = 12'h41D;
        15'h241A: data = 12'h407;
        15'h241B: data = 12'h3F7;
        15'h241C: data = 12'h3EA;
        15'h241D: data = 12'h3D2;
        15'h241E: data = 12'h3C3;
        15'h241F: data = 12'h3B2;
        15'h2420: data = 12'h39C;
        15'h2421: data = 12'h393;
        15'h2422: data = 12'h377;
        15'h2423: data = 12'h364;
        15'h2424: data = 12'h351;
        15'h2425: data = 12'h33D;
        15'h2426: data = 12'h330;
        15'h2427: data = 12'h320;
        15'h2428: data = 12'h30C;
        15'h2429: data = 12'h300;
        15'h242A: data = 12'h2EE;
        15'h242B: data = 12'h2E1;
        15'h242C: data = 12'h2D0;
        15'h242D: data = 12'h2D1;
        15'h242E: data = 12'h2C5;
        15'h242F: data = 12'h2B9;
        15'h2430: data = 12'h2AD;
        15'h2431: data = 12'h29D;
        15'h2432: data = 12'h297;
        15'h2433: data = 12'h286;
        15'h2434: data = 12'h27B;
        15'h2435: data = 12'h26A;
        15'h2436: data = 12'h25B;
        15'h2437: data = 12'h24B;
        15'h2438: data = 12'h242;
        15'h2439: data = 12'h230;
        15'h243A: data = 12'h224;
        15'h243B: data = 12'h213;
        15'h243C: data = 12'h20D;
        15'h243D: data = 12'h208;
        15'h243E: data = 12'h205;
        15'h243F: data = 12'h1F9;
        15'h2440: data = 12'h1F4;
        15'h2441: data = 12'h1EF;
        15'h2442: data = 12'h1EA;
        15'h2443: data = 12'h1E4;
        15'h2444: data = 12'h1D7;
        15'h2445: data = 12'h1C9;
        15'h2446: data = 12'h1C2;
        15'h2447: data = 12'h1B7;
        15'h2448: data = 12'h1B0;
        15'h2449: data = 12'h1A3;
        15'h244A: data = 12'h19A;
        15'h244B: data = 12'h190;
        15'h244C: data = 12'h194;
        15'h244D: data = 12'h18D;
        15'h244E: data = 12'h188;
        15'h244F: data = 12'h18C;
        15'h2450: data = 12'h18B;
        15'h2451: data = 12'h188;
        15'h2452: data = 12'h188;
        15'h2453: data = 12'h181;
        15'h2454: data = 12'h17D;
        15'h2455: data = 12'h175;
        15'h2456: data = 12'h173;
        15'h2457: data = 12'h170;
        15'h2458: data = 12'h164;
        15'h2459: data = 12'h15F;
        15'h245A: data = 12'h15F;
        15'h245B: data = 12'h15C;
        15'h245C: data = 12'h158;
        15'h245D: data = 12'h159;
        15'h245E: data = 12'h15A;
        15'h245F: data = 12'h161;
        15'h2460: data = 12'h164;
        15'h2461: data = 12'h164;
        15'h2462: data = 12'h16A;
        15'h2463: data = 12'h16D;
        15'h2464: data = 12'h16D;
        15'h2465: data = 12'h16B;
        15'h2466: data = 12'h16C;
        15'h2467: data = 12'h166;
        15'h2468: data = 12'h169;
        15'h2469: data = 12'h168;
        15'h246A: data = 12'h16B;
        15'h246B: data = 12'h16A;
        15'h246C: data = 12'h16B;
        15'h246D: data = 12'h178;
        15'h246E: data = 12'h180;
        15'h246F: data = 12'h187;
        15'h2470: data = 12'h18F;
        15'h2471: data = 12'h191;
        15'h2472: data = 12'h19D;
        15'h2473: data = 12'h1A3;
        15'h2474: data = 12'h1AD;
        15'h2475: data = 12'h1B0;
        15'h2476: data = 12'h1B2;
        15'h2477: data = 12'h1B5;
        15'h2478: data = 12'h1B9;
        15'h2479: data = 12'h1BC;
        15'h247A: data = 12'h1C5;
        15'h247B: data = 12'h1C8;
        15'h247C: data = 12'h1D0;
        15'h247D: data = 12'h1DA;
        15'h247E: data = 12'h1E3;
        15'h247F: data = 12'h1F0;
        15'h2480: data = 12'h200;
        15'h2481: data = 12'h20B;
        15'h2482: data = 12'h21B;
        15'h2483: data = 12'h221;
        15'h2484: data = 12'h22D;
        15'h2485: data = 12'h23A;
        15'h2486: data = 12'h248;
        15'h2487: data = 12'h24E;
        15'h2488: data = 12'h259;
        15'h2489: data = 12'h25D;
        15'h248A: data = 12'h26C;
        15'h248B: data = 12'h272;
        15'h248C: data = 12'h27A;
        15'h248D: data = 12'h283;
        15'h248E: data = 12'h291;
        15'h248F: data = 12'h2A0;
        15'h2490: data = 12'h2B7;
        15'h2491: data = 12'h2C3;
        15'h2492: data = 12'h2D4;
        15'h2493: data = 12'h2DE;
        15'h2494: data = 12'h2F5;
        15'h2495: data = 12'h307;
        15'h2496: data = 12'h318;
        15'h2497: data = 12'h328;
        15'h2498: data = 12'h338;
        15'h2499: data = 12'h343;
        15'h249A: data = 12'h355;
        15'h249B: data = 12'h360;
        15'h249C: data = 12'h36F;
        15'h249D: data = 12'h37D;
        15'h249E: data = 12'h392;
        15'h249F: data = 12'h396;
        15'h24A0: data = 12'h3A9;
        15'h24A1: data = 12'h3B9;
        15'h24A2: data = 12'h3C8;
        15'h24A3: data = 12'h3DB;
        15'h24A4: data = 12'h3EE;
        15'h24A5: data = 12'h3FE;
        15'h24A6: data = 12'h418;
        15'h24A7: data = 12'h42B;
        15'h24A8: data = 12'h443;
        15'h24A9: data = 12'h45A;
        15'h24AA: data = 12'h469;
        15'h24AB: data = 12'h483;
        15'h24AC: data = 12'h492;
        15'h24AD: data = 12'h4AA;
        15'h24AE: data = 12'h4B7;
        15'h24AF: data = 12'h4CF;
        15'h24B0: data = 12'h4E1;
        15'h24B1: data = 12'h4F7;
        15'h24B2: data = 12'h508;
        15'h24B3: data = 12'h51A;
        15'h24B4: data = 12'h52A;
        15'h24B5: data = 12'h53C;
        15'h24B6: data = 12'h553;
        15'h24B7: data = 12'h563;
        15'h24B8: data = 12'h577;
        15'h24B9: data = 12'h58C;
        15'h24BA: data = 12'h5A4;
        15'h24BB: data = 12'h5B6;
        15'h24BC: data = 12'h5CA;
        15'h24BD: data = 12'h5E5;
        15'h24BE: data = 12'h5FE;
        15'h24BF: data = 12'h61A;
        15'h24C0: data = 12'h62E;
        15'h24C1: data = 12'h647;
        15'h24C2: data = 12'h660;
        15'h24C3: data = 12'h677;
        15'h24C4: data = 12'h693;
        15'h24C5: data = 12'h6A5;
        15'h24C6: data = 12'h6B8;
        15'h24C7: data = 12'h6D0;
        15'h24C8: data = 12'h6E4;
        15'h24C9: data = 12'h6F5;
        15'h24CA: data = 12'h70B;
        15'h24CB: data = 12'h721;
        15'h24CC: data = 12'h736;
        15'h24CD: data = 12'h746;
        15'h24CE: data = 12'h75D;
        15'h24CF: data = 12'h773;
        15'h24D0: data = 12'h78E;
        15'h24D1: data = 12'h79F;
        15'h24D2: data = 12'h7B9;
        15'h24D3: data = 12'h7D7;
        15'h24D4: data = 12'h7EE;
        15'h24D5: data = 12'h804;
        15'h24D6: data = 12'h071;
        15'h24D7: data = 12'h08D;
        15'h24D8: data = 12'h0A1;
        15'h24D9: data = 12'h0B6;
        15'h24DA: data = 12'h0D4;
        15'h24DB: data = 12'h0E9;
        15'h24DC: data = 12'h100;
        15'h24DD: data = 12'h117;
        15'h24DE: data = 12'h12D;
        15'h24DF: data = 12'h144;
        15'h24E0: data = 12'h158;
        15'h24E1: data = 12'h16C;
        15'h24E2: data = 12'h181;
        15'h24E3: data = 12'h19C;
        15'h24E4: data = 12'h1B1;
        15'h24E5: data = 12'h1C0;
        15'h24E6: data = 12'h1D8;
        15'h24E7: data = 12'h1EF;
        15'h24E8: data = 12'h206;
        15'h24E9: data = 12'h218;
        15'h24EA: data = 12'h235;
        15'h24EB: data = 12'h24C;
        15'h24EC: data = 12'h262;
        15'h24ED: data = 12'h277;
        15'h24EE: data = 12'h28C;
        15'h24EF: data = 12'h2A8;
        15'h24F0: data = 12'h2C1;
        15'h24F1: data = 12'h2D7;
        15'h24F2: data = 12'h2F2;
        15'h24F3: data = 12'h309;
        15'h24F4: data = 12'h323;
        15'h24F5: data = 12'h33A;
        15'h24F6: data = 12'h34E;
        15'h24F7: data = 12'h369;
        15'h24F8: data = 12'h37C;
        15'h24F9: data = 12'h39E;
        15'h24FA: data = 12'h3AE;
        15'h24FB: data = 12'h3C6;
        15'h24FC: data = 12'h3DC;
        15'h24FD: data = 12'h3F3;
        15'h24FE: data = 12'h3FF;
        15'h24FF: data = 12'h418;
        15'h2500: data = 12'h42E;
        15'h2501: data = 12'h446;
        15'h2502: data = 12'h456;
        15'h2503: data = 12'h469;
        15'h2504: data = 12'h47C;
        15'h2505: data = 12'h496;
        15'h2506: data = 12'h4A7;
        15'h2507: data = 12'h4BA;
        15'h2508: data = 12'h4C9;
        15'h2509: data = 12'h4DB;
        15'h250A: data = 12'h4F0;
        15'h250B: data = 12'h507;
        15'h250C: data = 12'h513;
        15'h250D: data = 12'h527;
        15'h250E: data = 12'h53A;
        15'h250F: data = 12'h548;
        15'h2510: data = 12'h55E;
        15'h2511: data = 12'h56C;
        15'h2512: data = 12'h584;
        15'h2513: data = 12'h594;
        15'h2514: data = 12'h5A7;
        15'h2515: data = 12'h5BC;
        15'h2516: data = 12'h5C7;
        15'h2517: data = 12'h5D6;
        15'h2518: data = 12'h5F1;
        15'h2519: data = 12'h5FE;
        15'h251A: data = 12'h60E;
        15'h251B: data = 12'h61D;
        15'h251C: data = 12'h62F;
        15'h251D: data = 12'h63E;
        15'h251E: data = 12'h654;
        15'h251F: data = 12'h665;
        15'h2520: data = 12'h676;
        15'h2521: data = 12'h685;
        15'h2522: data = 12'h696;
        15'h2523: data = 12'h6A6;
        15'h2524: data = 12'h6B6;
        15'h2525: data = 12'h6C5;
        15'h2526: data = 12'h6D6;
        15'h2527: data = 12'h6DE;
        15'h2528: data = 12'h6EF;
        15'h2529: data = 12'h6FC;
        15'h252A: data = 12'h70C;
        15'h252B: data = 12'h718;
        15'h252C: data = 12'h725;
        15'h252D: data = 12'h736;
        15'h252E: data = 12'h73B;
        15'h252F: data = 12'h747;
        15'h2530: data = 12'h74F;
        15'h2531: data = 12'h760;
        15'h2532: data = 12'h767;
        15'h2533: data = 12'h776;
        15'h2534: data = 12'h77F;
        15'h2535: data = 12'h78E;
        15'h2536: data = 12'h799;
        15'h2537: data = 12'h79D;
        15'h2538: data = 12'h7A4;
        15'h2539: data = 12'h7AF;
        15'h253A: data = 12'h7B9;
        15'h253B: data = 12'h7BF;
        15'h253C: data = 12'h7C5;
        15'h253D: data = 12'h7CD;
        15'h253E: data = 12'h7D4;
        15'h253F: data = 12'h7DA;
        15'h2540: data = 12'h7E6;
        15'h2541: data = 12'h7EA;
        15'h2542: data = 12'h7F0;
        15'h2543: data = 12'h7FA;
        15'h2544: data = 12'h7FD;
        15'h2545: data = 12'h7FF;
        15'h2546: data = 12'h801;
        15'h2547: data = 12'h075;
        15'h2548: data = 12'h089;
        15'h2549: data = 12'h08A;
        15'h254A: data = 12'h097;
        15'h254B: data = 12'h098;
        15'h254C: data = 12'h099;
        15'h254D: data = 12'h0A4;
        15'h254E: data = 12'h0A0;
        15'h254F: data = 12'h0AD;
        15'h2550: data = 12'h0AB;
        15'h2551: data = 12'h0AE;
        15'h2552: data = 12'h0B8;
        15'h2553: data = 12'h0B9;
        15'h2554: data = 12'h0BD;
        15'h2555: data = 12'h0BD;
        15'h2556: data = 12'h0C8;
        15'h2557: data = 12'h0CD;
        15'h2558: data = 12'h0CE;
        15'h2559: data = 12'h0D2;
        15'h255A: data = 12'h0D4;
        15'h255B: data = 12'h0D7;
        15'h255C: data = 12'h0D7;
        15'h255D: data = 12'h0CE;
        15'h255E: data = 12'h0CF;
        15'h255F: data = 12'h0CA;
        15'h2560: data = 12'h0C7;
        15'h2561: data = 12'h0C5;
        15'h2562: data = 12'h0B8;
        15'h2563: data = 12'h0B6;
        15'h2564: data = 12'h0AF;
        15'h2565: data = 12'h0AF;
        15'h2566: data = 12'h0A8;
        15'h2567: data = 12'h0AB;
        15'h2568: data = 12'h0AF;
        15'h2569: data = 12'h0B2;
        15'h256A: data = 12'h0AD;
        15'h256B: data = 12'h0A4;
        15'h256C: data = 12'h0A3;
        15'h256D: data = 12'h098;
        15'h256E: data = 12'h08A;
        15'h256F: data = 12'h07D;
        15'h2570: data = 12'h071;
        15'h2571: data = 12'h075;
        15'h2572: data = 12'h073;
        15'h2573: data = 12'h070;
        15'h2574: data = 12'h06D;
        15'h2575: data = 12'h068;
        15'h2576: data = 12'h061;
        15'h2577: data = 12'h058;
        15'h2578: data = 12'h043;
        15'h2579: data = 12'h7BC;
        15'h257A: data = 12'h7B0;
        15'h257B: data = 12'h7AB;
        15'h257C: data = 12'h7A7;
        15'h257D: data = 12'h79E;
        15'h257E: data = 12'h796;
        15'h257F: data = 12'h78C;
        15'h2580: data = 12'h77B;
        15'h2581: data = 12'h76B;
        15'h2582: data = 12'h752;
        15'h2583: data = 12'h742;
        15'h2584: data = 12'h736;
        15'h2585: data = 12'h72F;
        15'h2586: data = 12'h727;
        15'h2587: data = 12'h722;
        15'h2588: data = 12'h718;
        15'h2589: data = 12'h70A;
        15'h258A: data = 12'h6F8;
        15'h258B: data = 12'h6E9;
        15'h258C: data = 12'h6D9;
        15'h258D: data = 12'h6C0;
        15'h258E: data = 12'h6B2;
        15'h258F: data = 12'h6A5;
        15'h2590: data = 12'h697;
        15'h2591: data = 12'h690;
        15'h2592: data = 12'h682;
        15'h2593: data = 12'h67A;
        15'h2594: data = 12'h668;
        15'h2595: data = 12'h65B;
        15'h2596: data = 12'h646;
        15'h2597: data = 12'h633;
        15'h2598: data = 12'h626;
        15'h2599: data = 12'h60A;
        15'h259A: data = 12'h5F7;
        15'h259B: data = 12'h5E3;
        15'h259C: data = 12'h5CD;
        15'h259D: data = 12'h5BF;
        15'h259E: data = 12'h5B3;
        15'h259F: data = 12'h5A7;
        15'h25A0: data = 12'h593;
        15'h25A1: data = 12'h589;
        15'h25A2: data = 12'h576;
        15'h25A3: data = 12'h569;
        15'h25A4: data = 12'h559;
        15'h25A5: data = 12'h543;
        15'h25A6: data = 12'h52C;
        15'h25A7: data = 12'h51A;
        15'h25A8: data = 12'h503;
        15'h25A9: data = 12'h4ED;
        15'h25AA: data = 12'h4D5;
        15'h25AB: data = 12'h4BF;
        15'h25AC: data = 12'h4AC;
        15'h25AD: data = 12'h495;
        15'h25AE: data = 12'h47C;
        15'h25AF: data = 12'h46A;
        15'h25B0: data = 12'h44F;
        15'h25B1: data = 12'h441;
        15'h25B2: data = 12'h42D;
        15'h25B3: data = 12'h416;
        15'h25B4: data = 12'h400;
        15'h25B5: data = 12'h3EA;
        15'h25B6: data = 12'h3D8;
        15'h25B7: data = 12'h3C3;
        15'h25B8: data = 12'h3B0;
        15'h25B9: data = 12'h397;
        15'h25BA: data = 12'h388;
        15'h25BB: data = 12'h370;
        15'h25BC: data = 12'h35F;
        15'h25BD: data = 12'h345;
        15'h25BE: data = 12'h336;
        15'h25BF: data = 12'h31C;
        15'h25C0: data = 12'h305;
        15'h25C1: data = 12'h2EF;
        15'h25C2: data = 12'h2DB;
        15'h25C3: data = 12'h2C9;
        15'h25C4: data = 12'h2AE;
        15'h25C5: data = 12'h292;
        15'h25C6: data = 12'h281;
        15'h25C7: data = 12'h268;
        15'h25C8: data = 12'h24F;
        15'h25C9: data = 12'h238;
        15'h25CA: data = 12'h21F;
        15'h25CB: data = 12'h20B;
        15'h25CC: data = 12'h1F6;
        15'h25CD: data = 12'h1D9;
        15'h25CE: data = 12'h1C1;
        15'h25CF: data = 12'h1AA;
        15'h25D0: data = 12'h194;
        15'h25D1: data = 12'h17C;
        15'h25D2: data = 12'h167;
        15'h25D3: data = 12'h14E;
        15'h25D4: data = 12'h137;
        15'h25D5: data = 12'h11F;
        15'h25D6: data = 12'h107;
        15'h25D7: data = 12'h0F3;
        15'h25D8: data = 12'h0DA;
        15'h25D9: data = 12'h0BE;
        15'h25DA: data = 12'h0A4;
        15'h25DB: data = 12'h08F;
        15'h25DC: data = 12'h080;
        15'h25DD: data = 12'h064;
        15'h25DE: data = 12'h04E;
        15'h25DF: data = 12'h7DD;
        15'h25E0: data = 12'h7CF;
        15'h25E1: data = 12'h7B9;
        15'h25E2: data = 12'h7A3;
        15'h25E3: data = 12'h78C;
        15'h25E4: data = 12'h776;
        15'h25E5: data = 12'h75B;
        15'h25E6: data = 12'h749;
        15'h25E7: data = 12'h734;
        15'h25E8: data = 12'h71A;
        15'h25E9: data = 12'h704;
        15'h25EA: data = 12'h6EC;
        15'h25EB: data = 12'h6D6;
        15'h25EC: data = 12'h6C3;
        15'h25ED: data = 12'h6AC;
        15'h25EE: data = 12'h697;
        15'h25EF: data = 12'h681;
        15'h25F0: data = 12'h667;
        15'h25F1: data = 12'h655;
        15'h25F2: data = 12'h638;
        15'h25F3: data = 12'h627;
        15'h25F4: data = 12'h613;
        15'h25F5: data = 12'h5F8;
        15'h25F6: data = 12'h5DF;
        15'h25F7: data = 12'h5CD;
        15'h25F8: data = 12'h5B6;
        15'h25F9: data = 12'h59E;
        15'h25FA: data = 12'h585;
        15'h25FB: data = 12'h56E;
        15'h25FC: data = 12'h55B;
        15'h25FD: data = 12'h546;
        15'h25FE: data = 12'h530;
        15'h25FF: data = 12'h51A;
        15'h2600: data = 12'h50A;
        15'h2601: data = 12'h4F3;
        15'h2602: data = 12'h4DC;
        15'h2603: data = 12'h4CC;
        15'h2604: data = 12'h4B9;
        15'h2605: data = 12'h4A5;
        15'h2606: data = 12'h492;
        15'h2607: data = 12'h47E;
        15'h2608: data = 12'h46E;
        15'h2609: data = 12'h45B;
        15'h260A: data = 12'h44D;
        15'h260B: data = 12'h441;
        15'h260C: data = 12'h42D;
        15'h260D: data = 12'h41B;
        15'h260E: data = 12'h407;
        15'h260F: data = 12'h3FB;
        15'h2610: data = 12'h3EA;
        15'h2611: data = 12'h3D3;
        15'h2612: data = 12'h3C1;
        15'h2613: data = 12'h3AF;
        15'h2614: data = 12'h39B;
        15'h2615: data = 12'h38E;
        15'h2616: data = 12'h376;
        15'h2617: data = 12'h361;
        15'h2618: data = 12'h350;
        15'h2619: data = 12'h33D;
        15'h261A: data = 12'h32D;
        15'h261B: data = 12'h31D;
        15'h261C: data = 12'h30E;
        15'h261D: data = 12'h2FF;
        15'h261E: data = 12'h2F2;
        15'h261F: data = 12'h2E3;
        15'h2620: data = 12'h2DA;
        15'h2621: data = 12'h2D5;
        15'h2622: data = 12'h2C8;
        15'h2623: data = 12'h2BC;
        15'h2624: data = 12'h2AD;
        15'h2625: data = 12'h2A3;
        15'h2626: data = 12'h292;
        15'h2627: data = 12'h284;
        15'h2628: data = 12'h279;
        15'h2629: data = 12'h264;
        15'h262A: data = 12'h25B;
        15'h262B: data = 12'h246;
        15'h262C: data = 12'h23D;
        15'h262D: data = 12'h22B;
        15'h262E: data = 12'h221;
        15'h262F: data = 12'h217;
        15'h2630: data = 12'h212;
        15'h2631: data = 12'h20D;
        15'h2632: data = 12'h20A;
        15'h2633: data = 12'h1FD;
        15'h2634: data = 12'h1FB;
        15'h2635: data = 12'h1F3;
        15'h2636: data = 12'h1EC;
        15'h2637: data = 12'h1E4;
        15'h2638: data = 12'h1D3;
        15'h2639: data = 12'h1C9;
        15'h263A: data = 12'h1BE;
        15'h263B: data = 12'h1B8;
        15'h263C: data = 12'h1AD;
        15'h263D: data = 12'h1A3;
        15'h263E: data = 12'h19A;
        15'h263F: data = 12'h195;
        15'h2640: data = 12'h194;
        15'h2641: data = 12'h18F;
        15'h2642: data = 12'h18F;
        15'h2643: data = 12'h18D;
        15'h2644: data = 12'h18D;
        15'h2645: data = 12'h188;
        15'h2646: data = 12'h187;
        15'h2647: data = 12'h180;
        15'h2648: data = 12'h179;
        15'h2649: data = 12'h172;
        15'h264A: data = 12'h16D;
        15'h264B: data = 12'h169;
        15'h264C: data = 12'h15D;
        15'h264D: data = 12'h15B;
        15'h264E: data = 12'h15F;
        15'h264F: data = 12'h15C;
        15'h2650: data = 12'h158;
        15'h2651: data = 12'h15F;
        15'h2652: data = 12'h163;
        15'h2653: data = 12'h168;
        15'h2654: data = 12'h168;
        15'h2655: data = 12'h169;
        15'h2656: data = 12'h169;
        15'h2657: data = 12'h170;
        15'h2658: data = 12'h16D;
        15'h2659: data = 12'h16D;
        15'h265A: data = 12'h168;
        15'h265B: data = 12'h165;
        15'h265C: data = 12'h16A;
        15'h265D: data = 12'h166;
        15'h265E: data = 12'h16A;
        15'h265F: data = 12'h16E;
        15'h2660: data = 12'h16F;
        15'h2661: data = 12'h17A;
        15'h2662: data = 12'h186;
        15'h2663: data = 12'h188;
        15'h2664: data = 12'h197;
        15'h2665: data = 12'h197;
        15'h2666: data = 12'h19E;
        15'h2667: data = 12'h1A4;
        15'h2668: data = 12'h1AF;
        15'h2669: data = 12'h1B1;
        15'h266A: data = 12'h1AD;
        15'h266B: data = 12'h1B4;
        15'h266C: data = 12'h1B6;
        15'h266D: data = 12'h1C0;
        15'h266E: data = 12'h1C2;
        15'h266F: data = 12'h1C9;
        15'h2670: data = 12'h1D0;
        15'h2671: data = 12'h1DB;
        15'h2672: data = 12'h1E5;
        15'h2673: data = 12'h1F7;
        15'h2674: data = 12'h200;
        15'h2675: data = 12'h20E;
        15'h2676: data = 12'h21C;
        15'h2677: data = 12'h222;
        15'h2678: data = 12'h232;
        15'h2679: data = 12'h239;
        15'h267A: data = 12'h247;
        15'h267B: data = 12'h24C;
        15'h267C: data = 12'h25A;
        15'h267D: data = 12'h25E;
        15'h267E: data = 12'h26A;
        15'h267F: data = 12'h26E;
        15'h2680: data = 12'h27C;
        15'h2681: data = 12'h286;
        15'h2682: data = 12'h293;
        15'h2683: data = 12'h2A2;
        15'h2684: data = 12'h2B5;
        15'h2685: data = 12'h2C5;
        15'h2686: data = 12'h2D9;
        15'h2687: data = 12'h2E2;
        15'h2688: data = 12'h2F8;
        15'h2689: data = 12'h309;
        15'h268A: data = 12'h316;
        15'h268B: data = 12'h327;
        15'h268C: data = 12'h337;
        15'h268D: data = 12'h344;
        15'h268E: data = 12'h355;
        15'h268F: data = 12'h362;
        15'h2690: data = 12'h36F;
        15'h2691: data = 12'h37D;
        15'h2692: data = 12'h38E;
        15'h2693: data = 12'h395;
        15'h2694: data = 12'h3AB;
        15'h2695: data = 12'h3B7;
        15'h2696: data = 12'h3C7;
        15'h2697: data = 12'h3DE;
        15'h2698: data = 12'h3F0;
        15'h2699: data = 12'h402;
        15'h269A: data = 12'h41C;
        15'h269B: data = 12'h42F;
        15'h269C: data = 12'h446;
        15'h269D: data = 12'h458;
        15'h269E: data = 12'h46F;
        15'h269F: data = 12'h483;
        15'h26A0: data = 12'h494;
        15'h26A1: data = 12'h4AD;
        15'h26A2: data = 12'h4B8;
        15'h26A3: data = 12'h4CF;
        15'h26A4: data = 12'h4E5;
        15'h26A5: data = 12'h4F4;
        15'h26A6: data = 12'h506;
        15'h26A7: data = 12'h515;
        15'h26A8: data = 12'h528;
        15'h26A9: data = 12'h53D;
        15'h26AA: data = 12'h555;
        15'h26AB: data = 12'h567;
        15'h26AC: data = 12'h578;
        15'h26AD: data = 12'h591;
        15'h26AE: data = 12'h5A1;
        15'h26AF: data = 12'h5B9;
        15'h26B0: data = 12'h5CF;
        15'h26B1: data = 12'h5EC;
        15'h26B2: data = 12'h603;
        15'h26B3: data = 12'h620;
        15'h26B4: data = 12'h634;
        15'h26B5: data = 12'h64E;
        15'h26B6: data = 12'h665;
        15'h26B7: data = 12'h67B;
        15'h26B8: data = 12'h691;
        15'h26B9: data = 12'h6A1;
        15'h26BA: data = 12'h6B5;
        15'h26BB: data = 12'h6CC;
        15'h26BC: data = 12'h6DF;
        15'h26BD: data = 12'h6F5;
        15'h26BE: data = 12'h709;
        15'h26BF: data = 12'h71D;
        15'h26C0: data = 12'h735;
        15'h26C1: data = 12'h743;
        15'h26C2: data = 12'h75D;
        15'h26C3: data = 12'h774;
        15'h26C4: data = 12'h791;
        15'h26C5: data = 12'h7A4;
        15'h26C6: data = 12'h7BA;
        15'h26C7: data = 12'h7D8;
        15'h26C8: data = 12'h7F0;
        15'h26C9: data = 12'h806;
        15'h26CA: data = 12'h073;
        15'h26CB: data = 12'h08F;
        15'h26CC: data = 12'h0A2;
        15'h26CD: data = 12'h0B8;
        15'h26CE: data = 12'h0D2;
        15'h26CF: data = 12'h0EA;
        15'h26D0: data = 12'h101;
        15'h26D1: data = 12'h116;
        15'h26D2: data = 12'h12B;
        15'h26D3: data = 12'h147;
        15'h26D4: data = 12'h155;
        15'h26D5: data = 12'h16B;
        15'h26D6: data = 12'h180;
        15'h26D7: data = 12'h198;
        15'h26D8: data = 12'h1AD;
        15'h26D9: data = 12'h1BE;
        15'h26DA: data = 12'h1D7;
        15'h26DB: data = 12'h1EF;
        15'h26DC: data = 12'h207;
        15'h26DD: data = 12'h21B;
        15'h26DE: data = 12'h232;
        15'h26DF: data = 12'h249;
        15'h26E0: data = 12'h263;
        15'h26E1: data = 12'h27A;
        15'h26E2: data = 12'h290;
        15'h26E3: data = 12'h2AB;
        15'h26E4: data = 12'h2C3;
        15'h26E5: data = 12'h2DB;
        15'h26E6: data = 12'h2F3;
        15'h26E7: data = 12'h30C;
        15'h26E8: data = 12'h329;
        15'h26E9: data = 12'h33B;
        15'h26EA: data = 12'h353;
        15'h26EB: data = 12'h36C;
        15'h26EC: data = 12'h382;
        15'h26ED: data = 12'h39C;
        15'h26EE: data = 12'h3AB;
        15'h26EF: data = 12'h3C3;
        15'h26F0: data = 12'h3DD;
        15'h26F1: data = 12'h3F0;
        15'h26F2: data = 12'h3FE;
        15'h26F3: data = 12'h416;
        15'h26F4: data = 12'h42C;
        15'h26F5: data = 12'h442;
        15'h26F6: data = 12'h453;
        15'h26F7: data = 12'h467;
        15'h26F8: data = 12'h47E;
        15'h26F9: data = 12'h492;
        15'h26FA: data = 12'h4A5;
        15'h26FB: data = 12'h4B7;
        15'h26FC: data = 12'h4C4;
        15'h26FD: data = 12'h4D7;
        15'h26FE: data = 12'h4EF;
        15'h26FF: data = 12'h505;
        15'h2700: data = 12'h511;
        15'h2701: data = 12'h525;
        15'h2702: data = 12'h53C;
        15'h2703: data = 12'h548;
        15'h2704: data = 12'h55C;
        15'h2705: data = 12'h571;
        15'h2706: data = 12'h584;
        15'h2707: data = 12'h593;
        15'h2708: data = 12'h5A4;
        15'h2709: data = 12'h5B8;
        15'h270A: data = 12'h5C3;
        15'h270B: data = 12'h5D7;
        15'h270C: data = 12'h5EE;
        15'h270D: data = 12'h5FE;
        15'h270E: data = 12'h60F;
        15'h270F: data = 12'h61E;
        15'h2710: data = 12'h630;
        15'h2711: data = 12'h640;
        15'h2712: data = 12'h655;
        15'h2713: data = 12'h666;
        15'h2714: data = 12'h679;
        15'h2715: data = 12'h689;
        15'h2716: data = 12'h698;
        15'h2717: data = 12'h6A7;
        15'h2718: data = 12'h6B4;
        15'h2719: data = 12'h6C5;
        15'h271A: data = 12'h6D4;
        15'h271B: data = 12'h6DF;
        15'h271C: data = 12'h6EF;
        15'h271D: data = 12'h6FE;
        15'h271E: data = 12'h70A;
        15'h271F: data = 12'h714;
        15'h2720: data = 12'h727;
        15'h2721: data = 12'h736;
        15'h2722: data = 12'h739;
        15'h2723: data = 12'h749;
        15'h2724: data = 12'h751;
        15'h2725: data = 12'h75F;
        15'h2726: data = 12'h766;
        15'h2727: data = 12'h775;
        15'h2728: data = 12'h77C;
        15'h2729: data = 12'h78F;
        15'h272A: data = 12'h794;
        15'h272B: data = 12'h79D;
        15'h272C: data = 12'h7A3;
        15'h272D: data = 12'h7B1;
        15'h272E: data = 12'h7B8;
        15'h272F: data = 12'h7BE;
        15'h2730: data = 12'h7C3;
        15'h2731: data = 12'h7CE;
        15'h2732: data = 12'h7D1;
        15'h2733: data = 12'h7D9;
        15'h2734: data = 12'h7E5;
        15'h2735: data = 12'h7E5;
        15'h2736: data = 12'h7ED;
        15'h2737: data = 12'h7F2;
        15'h2738: data = 12'h7FC;
        15'h2739: data = 12'h7FD;
        15'h273A: data = 12'h800;
        15'h273B: data = 12'h80A;
        15'h273C: data = 12'h077;
        15'h273D: data = 12'h089;
        15'h273E: data = 12'h093;
        15'h273F: data = 12'h096;
        15'h2740: data = 12'h094;
        15'h2741: data = 12'h0A1;
        15'h2742: data = 12'h0A3;
        15'h2743: data = 12'h0AB;
        15'h2744: data = 12'h0AC;
        15'h2745: data = 12'h0AE;
        15'h2746: data = 12'h0B7;
        15'h2747: data = 12'h0B9;
        15'h2748: data = 12'h0BF;
        15'h2749: data = 12'h0BF;
        15'h274A: data = 12'h0C8;
        15'h274B: data = 12'h0CF;
        15'h274C: data = 12'h0D1;
        15'h274D: data = 12'h0D3;
        15'h274E: data = 12'h0D3;
        15'h274F: data = 12'h0D6;
        15'h2750: data = 12'h0D5;
        15'h2751: data = 12'h0CD;
        15'h2752: data = 12'h0CC;
        15'h2753: data = 12'h0CA;
        15'h2754: data = 12'h0C9;
        15'h2755: data = 12'h0C3;
        15'h2756: data = 12'h0B9;
        15'h2757: data = 12'h0B7;
        15'h2758: data = 12'h0AD;
        15'h2759: data = 12'h0AE;
        15'h275A: data = 12'h0A8;
        15'h275B: data = 12'h0AF;
        15'h275C: data = 12'h0B1;
        15'h275D: data = 12'h0B5;
        15'h275E: data = 12'h0AE;
        15'h275F: data = 12'h0A6;
        15'h2760: data = 12'h0A3;
        15'h2761: data = 12'h09D;
        15'h2762: data = 12'h08E;
        15'h2763: data = 12'h084;
        15'h2764: data = 12'h075;
        15'h2765: data = 12'h077;
        15'h2766: data = 12'h071;
        15'h2767: data = 12'h06D;
        15'h2768: data = 12'h06F;
        15'h2769: data = 12'h069;
        15'h276A: data = 12'h061;
        15'h276B: data = 12'h059;
        15'h276C: data = 12'h048;
        15'h276D: data = 12'h032;
        15'h276E: data = 12'h7B7;
        15'h276F: data = 12'h7AE;
        15'h2770: data = 12'h7A5;
        15'h2771: data = 12'h79E;
        15'h2772: data = 12'h799;
        15'h2773: data = 12'h791;
        15'h2774: data = 12'h781;
        15'h2775: data = 12'h771;
        15'h2776: data = 12'h75B;
        15'h2777: data = 12'h746;
        15'h2778: data = 12'h736;
        15'h2779: data = 12'h730;
        15'h277A: data = 12'h72C;
        15'h277B: data = 12'h720;
        15'h277C: data = 12'h718;
        15'h277D: data = 12'h711;
        15'h277E: data = 12'h6FD;
        15'h277F: data = 12'h6EA;
        15'h2780: data = 12'h6DE;
        15'h2781: data = 12'h6C7;
        15'h2782: data = 12'h6B5;
        15'h2783: data = 12'h6A9;
        15'h2784: data = 12'h695;
        15'h2785: data = 12'h68C;
        15'h2786: data = 12'h684;
        15'h2787: data = 12'h678;
        15'h2788: data = 12'h66A;
        15'h2789: data = 12'h65A;
        15'h278A: data = 12'h646;
        15'h278B: data = 12'h635;
        15'h278C: data = 12'h62B;
        15'h278D: data = 12'h609;
        15'h278E: data = 12'h5F6;
        15'h278F: data = 12'h5E5;
        15'h2790: data = 12'h5D0;
        15'h2791: data = 12'h5C1;
        15'h2792: data = 12'h5B4;
        15'h2793: data = 12'h5A9;
        15'h2794: data = 12'h595;
        15'h2795: data = 12'h589;
        15'h2796: data = 12'h579;
        15'h2797: data = 12'h567;
        15'h2798: data = 12'h55A;
        15'h2799: data = 12'h547;
        15'h279A: data = 12'h52C;
        15'h279B: data = 12'h51A;
        15'h279C: data = 12'h502;
        15'h279D: data = 12'h4F0;
        15'h279E: data = 12'h4D6;
        15'h279F: data = 12'h4C1;
        15'h27A0: data = 12'h4AC;
        15'h27A1: data = 12'h496;
        15'h27A2: data = 12'h480;
        15'h27A3: data = 12'h46C;
        15'h27A4: data = 12'h453;
        15'h27A5: data = 12'h440;
        15'h27A6: data = 12'h42C;
        15'h27A7: data = 12'h41A;
        15'h27A8: data = 12'h402;
        15'h27A9: data = 12'h3ED;
        15'h27AA: data = 12'h3DB;
        15'h27AB: data = 12'h3C8;
        15'h27AC: data = 12'h3B7;
        15'h27AD: data = 12'h39B;
        15'h27AE: data = 12'h38C;
        15'h27AF: data = 12'h376;
        15'h27B0: data = 12'h35E;
        15'h27B1: data = 12'h347;
        15'h27B2: data = 12'h331;
        15'h27B3: data = 12'h320;
        15'h27B4: data = 12'h308;
        15'h27B5: data = 12'h2F2;
        15'h27B6: data = 12'h2DC;
        15'h27B7: data = 12'h2C7;
        15'h27B8: data = 12'h2AD;
        15'h27B9: data = 12'h294;
        15'h27BA: data = 12'h283;
        15'h27BB: data = 12'h26C;
        15'h27BC: data = 12'h250;
        15'h27BD: data = 12'h23A;
        15'h27BE: data = 12'h21F;
        15'h27BF: data = 12'h209;
        15'h27C0: data = 12'h1F4;
        15'h27C1: data = 12'h1DB;
        15'h27C2: data = 12'h1C1;
        15'h27C3: data = 12'h1AC;
        15'h27C4: data = 12'h195;
        15'h27C5: data = 12'h181;
        15'h27C6: data = 12'h165;
        15'h27C7: data = 12'h14F;
        15'h27C8: data = 12'h137;
        15'h27C9: data = 12'h11F;
        15'h27CA: data = 12'h10B;
        15'h27CB: data = 12'h0F4;
        15'h27CC: data = 12'h0DF;
        15'h27CD: data = 12'h0C1;
        15'h27CE: data = 12'h0A9;
        15'h27CF: data = 12'h091;
        15'h27D0: data = 12'h07F;
        15'h27D1: data = 12'h064;
        15'h27D2: data = 12'h04A;
        15'h27D3: data = 12'h6BE;
        15'h27D4: data = 12'h7CD;
        15'h27D5: data = 12'h7B7;
        15'h27D6: data = 12'h7A2;
        15'h27D7: data = 12'h78B;
        15'h27D8: data = 12'h774;
        15'h27D9: data = 12'h75B;
        15'h27DA: data = 12'h74B;
        15'h27DB: data = 12'h735;
        15'h27DC: data = 12'h71D;
        15'h27DD: data = 12'h705;
        15'h27DE: data = 12'h6EC;
        15'h27DF: data = 12'h6D5;
        15'h27E0: data = 12'h6C0;
        15'h27E1: data = 12'h6A9;
        15'h27E2: data = 12'h693;
        15'h27E3: data = 12'h67E;
        15'h27E4: data = 12'h665;
        15'h27E5: data = 12'h651;
        15'h27E6: data = 12'h638;
        15'h27E7: data = 12'h624;
        15'h27E8: data = 12'h60E;
        15'h27E9: data = 12'h5F3;
        15'h27EA: data = 12'h5DB;
        15'h27EB: data = 12'h5C5;
        15'h27EC: data = 12'h5B5;
        15'h27ED: data = 12'h598;
        15'h27EE: data = 12'h582;
        15'h27EF: data = 12'h56C;
        15'h27F0: data = 12'h55A;
        15'h27F1: data = 12'h547;
        15'h27F2: data = 12'h531;
        15'h27F3: data = 12'h51A;
        15'h27F4: data = 12'h50A;
        15'h27F5: data = 12'h4F4;
        15'h27F6: data = 12'h4DF;
        15'h27F7: data = 12'h4D0;
        15'h27F8: data = 12'h4BC;
        15'h27F9: data = 12'h4AB;
        15'h27FA: data = 12'h498;
        15'h27FB: data = 12'h488;
        15'h27FC: data = 12'h475;
        15'h27FD: data = 12'h464;
        15'h27FE: data = 12'h454;
        15'h27FF: data = 12'h446;
        15'h2800: data = 12'h42F;
        15'h2801: data = 12'h41D;
        15'h2802: data = 12'h40A;
        15'h2803: data = 12'h3F8;
        15'h2804: data = 12'h3E9;
        15'h2805: data = 12'h3D2;
        15'h2806: data = 12'h3C2;
        15'h2807: data = 12'h3B0;
        15'h2808: data = 12'h39B;
        15'h2809: data = 12'h38E;
        15'h280A: data = 12'h373;
        15'h280B: data = 12'h35C;
        15'h280C: data = 12'h34F;
        15'h280D: data = 12'h33D;
        15'h280E: data = 12'h32C;
        15'h280F: data = 12'h31E;
        15'h2810: data = 12'h310;
        15'h2811: data = 12'h300;
        15'h2812: data = 12'h2F3;
        15'h2813: data = 12'h2E8;
        15'h2814: data = 12'h2DD;
        15'h2815: data = 12'h2D8;
        15'h2816: data = 12'h2CA;
        15'h2817: data = 12'h2BF;
        15'h2818: data = 12'h2AC;
        15'h2819: data = 12'h2A2;
        15'h281A: data = 12'h293;
        15'h281B: data = 12'h283;
        15'h281C: data = 12'h278;
        15'h281D: data = 12'h264;
        15'h281E: data = 12'h258;
        15'h281F: data = 12'h24A;
        15'h2820: data = 12'h240;
        15'h2821: data = 12'h22B;
        15'h2822: data = 12'h222;
        15'h2823: data = 12'h21A;
        15'h2824: data = 12'h214;
        15'h2825: data = 12'h212;
        15'h2826: data = 12'h20D;
        15'h2827: data = 12'h200;
        15'h2828: data = 12'h1FC;
        15'h2829: data = 12'h1F1;
        15'h282A: data = 12'h1ED;
        15'h282B: data = 12'h1E4;
        15'h282C: data = 12'h1D6;
        15'h282D: data = 12'h1C8;
        15'h282E: data = 12'h1BA;
        15'h282F: data = 12'h1B7;
        15'h2830: data = 12'h1AB;
        15'h2831: data = 12'h1A1;
        15'h2832: data = 12'h19B;
        15'h2833: data = 12'h195;
        15'h2834: data = 12'h193;
        15'h2835: data = 12'h193;
        15'h2836: data = 12'h18F;
        15'h2837: data = 12'h192;
        15'h2838: data = 12'h18F;
        15'h2839: data = 12'h188;
        15'h283A: data = 12'h186;
        15'h283B: data = 12'h17E;
        15'h283C: data = 12'h17E;
        15'h283D: data = 12'h171;
        15'h283E: data = 12'h16B;
        15'h283F: data = 12'h169;
        15'h2840: data = 12'h15D;
        15'h2841: data = 12'h15D;
        15'h2842: data = 12'h15C;
        15'h2843: data = 12'h15F;
        15'h2844: data = 12'h156;
        15'h2845: data = 12'h15D;
        15'h2846: data = 12'h163;
        15'h2847: data = 12'h166;
        15'h2848: data = 12'h168;
        15'h2849: data = 12'h166;
        15'h284A: data = 12'h167;
        15'h284B: data = 12'h171;
        15'h284C: data = 12'h16A;
        15'h284D: data = 12'h165;
        15'h284E: data = 12'h162;
        15'h284F: data = 12'h15F;
        15'h2850: data = 12'h164;
        15'h2851: data = 12'h163;
        15'h2852: data = 12'h16B;
        15'h2853: data = 12'h16C;
        15'h2854: data = 12'h16E;
        15'h2855: data = 12'h17D;
        15'h2856: data = 12'h188;
        15'h2857: data = 12'h18D;
        15'h2858: data = 12'h194;
        15'h2859: data = 12'h194;
        15'h285A: data = 12'h19C;
        15'h285B: data = 12'h1A0;
        15'h285C: data = 12'h1A9;
        15'h285D: data = 12'h1B0;
        15'h285E: data = 12'h1AA;
        15'h285F: data = 12'h1AD;
        15'h2860: data = 12'h1B5;
        15'h2861: data = 12'h1BA;
        15'h2862: data = 12'h1BF;
        15'h2863: data = 12'h1C9;
        15'h2864: data = 12'h1D0;
        15'h2865: data = 12'h1DA;
        15'h2866: data = 12'h1E7;
        15'h2867: data = 12'h1F8;
        15'h2868: data = 12'h207;
        15'h2869: data = 12'h20F;
        15'h286A: data = 12'h21D;
        15'h286B: data = 12'h222;
        15'h286C: data = 12'h22C;
        15'h286D: data = 12'h234;
        15'h286E: data = 12'h245;
        15'h286F: data = 12'h249;
        15'h2870: data = 12'h258;
        15'h2871: data = 12'h25A;
        15'h2872: data = 12'h267;
        15'h2873: data = 12'h26B;
        15'h2874: data = 12'h278;
        15'h2875: data = 12'h287;
        15'h2876: data = 12'h294;
        15'h2877: data = 12'h2A3;
        15'h2878: data = 12'h2B5;
        15'h2879: data = 12'h2C8;
        15'h287A: data = 12'h2D9;
        15'h287B: data = 12'h2E5;
        15'h287C: data = 12'h2F7;
        15'h287D: data = 12'h307;
        15'h287E: data = 12'h319;
        15'h287F: data = 12'h326;
        15'h2880: data = 12'h333;
        15'h2881: data = 12'h341;
        15'h2882: data = 12'h34E;
        15'h2883: data = 12'h35B;
        15'h2884: data = 12'h36A;
        15'h2885: data = 12'h375;
        15'h2886: data = 12'h389;
        15'h2887: data = 12'h38F;
        15'h2888: data = 12'h3A8;
        15'h2889: data = 12'h3B7;
        15'h288A: data = 12'h3C7;
        15'h288B: data = 12'h3E1;
        15'h288C: data = 12'h3F0;
        15'h288D: data = 12'h403;
        15'h288E: data = 12'h41D;
        15'h288F: data = 12'h432;
        15'h2890: data = 12'h44A;
        15'h2891: data = 12'h45A;
        15'h2892: data = 12'h46C;
        15'h2893: data = 12'h482;
        15'h2894: data = 12'h491;
        15'h2895: data = 12'h4A7;
        15'h2896: data = 12'h4B7;
        15'h2897: data = 12'h4CB;
        15'h2898: data = 12'h4DB;
        15'h2899: data = 12'h4EB;
        15'h289A: data = 12'h500;
        15'h289B: data = 12'h510;
        15'h289C: data = 12'h526;
        15'h289D: data = 12'h53A;
        15'h289E: data = 12'h550;
        15'h289F: data = 12'h564;
        15'h28A0: data = 12'h575;
        15'h28A1: data = 12'h58A;
        15'h28A2: data = 12'h5A6;
        15'h28A3: data = 12'h5C0;
        15'h28A4: data = 12'h5D4;
        15'h28A5: data = 12'h5EE;
        15'h28A6: data = 12'h606;
        15'h28A7: data = 12'h61F;
        15'h28A8: data = 12'h634;
        15'h28A9: data = 12'h64A;
        15'h28AA: data = 12'h660;
        15'h28AB: data = 12'h675;
        15'h28AC: data = 12'h691;
        15'h28AD: data = 12'h69D;
        15'h28AE: data = 12'h6B3;
        15'h28AF: data = 12'h6CA;
        15'h28B0: data = 12'h6DC;
        15'h28B1: data = 12'h6EE;
        15'h28B2: data = 12'h703;
        15'h28B3: data = 12'h714;
        15'h28B4: data = 12'h72F;
        15'h28B5: data = 12'h742;
        15'h28B6: data = 12'h757;
        15'h28B7: data = 12'h773;
        15'h28B8: data = 12'h790;
        15'h28B9: data = 12'h7A2;
        15'h28BA: data = 12'h7BD;
        15'h28BB: data = 12'h7DC;
        15'h28BC: data = 12'h7F3;
        15'h28BD: data = 12'h809;
        15'h28BE: data = 12'h078;
        15'h28BF: data = 12'h08C;
        15'h28C0: data = 12'h0A5;
        15'h28C1: data = 12'h0BA;
        15'h28C2: data = 12'h0D2;
        15'h28C3: data = 12'h0E7;
        15'h28C4: data = 12'h0FE;
        15'h28C5: data = 12'h10E;
        15'h28C6: data = 12'h124;
        15'h28C7: data = 12'h13F;
        15'h28C8: data = 12'h151;
        15'h28C9: data = 12'h162;
        15'h28CA: data = 12'h179;
        15'h28CB: data = 12'h18F;
        15'h28CC: data = 12'h1A8;
        15'h28CD: data = 12'h1B7;
        15'h28CE: data = 12'h1D3;
        15'h28CF: data = 12'h1E9;
        15'h28D0: data = 12'h205;
        15'h28D1: data = 12'h21A;
        15'h28D2: data = 12'h233;
        15'h28D3: data = 12'h24C;
        15'h28D4: data = 12'h264;
        15'h28D5: data = 12'h279;
        15'h28D6: data = 12'h292;
        15'h28D7: data = 12'h2AE;
        15'h28D8: data = 12'h2C7;
        15'h28D9: data = 12'h2DD;
        15'h28DA: data = 12'h2F9;
        15'h28DB: data = 12'h310;
        15'h28DC: data = 12'h32A;
        15'h28DD: data = 12'h33A;
        15'h28DE: data = 12'h351;
        15'h28DF: data = 12'h369;
        15'h28E0: data = 12'h37F;
        15'h28E1: data = 12'h398;
        15'h28E2: data = 12'h3AA;
        15'h28E3: data = 12'h3C2;
        15'h28E4: data = 12'h3D9;
        15'h28E5: data = 12'h3EC;
        15'h28E6: data = 12'h3FC;
        15'h28E7: data = 12'h411;
        15'h28E8: data = 12'h429;
        15'h28E9: data = 12'h43E;
        15'h28EA: data = 12'h44B;
        15'h28EB: data = 12'h45D;
        15'h28EC: data = 12'h475;
        15'h28ED: data = 12'h48A;
        15'h28EE: data = 12'h49F;
        15'h28EF: data = 12'h4B0;
        15'h28F0: data = 12'h4C1;
        15'h28F1: data = 12'h4D6;
        15'h28F2: data = 12'h4EB;
        15'h28F3: data = 12'h500;
        15'h28F4: data = 12'h50B;
        15'h28F5: data = 12'h523;
        15'h28F6: data = 12'h53B;
        15'h28F7: data = 12'h549;
        15'h28F8: data = 12'h55A;
        15'h28F9: data = 12'h56C;
        15'h28FA: data = 12'h583;
        15'h28FB: data = 12'h590;
        15'h28FC: data = 12'h5A8;
        15'h28FD: data = 12'h5BE;
        15'h28FE: data = 12'h5CC;
        15'h28FF: data = 12'h5DC;
        15'h2900: data = 12'h5F4;
        15'h2901: data = 12'h605;
        15'h2902: data = 12'h615;
        15'h2903: data = 12'h626;
        15'h2904: data = 12'h637;
        15'h2905: data = 12'h648;
        15'h2906: data = 12'h65C;
        15'h2907: data = 12'h669;
        15'h2908: data = 12'h67B;
        15'h2909: data = 12'h68A;
        15'h290A: data = 12'h69D;
        15'h290B: data = 12'h6AA;
        15'h290C: data = 12'h6BB;
        15'h290D: data = 12'h6C6;
        15'h290E: data = 12'h6D8;
        15'h290F: data = 12'h6E1;
        15'h2910: data = 12'h6F0;
        15'h2911: data = 12'h701;
        15'h2912: data = 12'h70C;
        15'h2913: data = 12'h715;
        15'h2914: data = 12'h726;
        15'h2915: data = 12'h733;
        15'h2916: data = 12'h73A;
        15'h2917: data = 12'h747;
        15'h2918: data = 12'h74E;
        15'h2919: data = 12'h75E;
        15'h291A: data = 12'h765;
        15'h291B: data = 12'h774;
        15'h291C: data = 12'h77D;
        15'h291D: data = 12'h789;
        15'h291E: data = 12'h791;
        15'h291F: data = 12'h79C;
        15'h2920: data = 12'h7A2;
        15'h2921: data = 12'h7AB;
        15'h2922: data = 12'h7B0;
        15'h2923: data = 12'h7B7;
        15'h2924: data = 12'h7C0;
        15'h2925: data = 12'h7C7;
        15'h2926: data = 12'h7CC;
        15'h2927: data = 12'h7D4;
        15'h2928: data = 12'h7DD;
        15'h2929: data = 12'h7E2;
        15'h292A: data = 12'h7EA;
        15'h292B: data = 12'h7F0;
        15'h292C: data = 12'h7F8;
        15'h292D: data = 12'h7FA;
        15'h292E: data = 12'h7FF;
        15'h292F: data = 12'h802;
        15'h2930: data = 12'h521;
        15'h2931: data = 12'h085;
        15'h2932: data = 12'h08F;
        15'h2933: data = 12'h093;
        15'h2934: data = 12'h092;
        15'h2935: data = 12'h09F;
        15'h2936: data = 12'h0A1;
        15'h2937: data = 12'h0AD;
        15'h2938: data = 12'h0AB;
        15'h2939: data = 12'h0B0;
        15'h293A: data = 12'h0B9;
        15'h293B: data = 12'h0B9;
        15'h293C: data = 12'h0BE;
        15'h293D: data = 12'h0C0;
        15'h293E: data = 12'h0CD;
        15'h293F: data = 12'h0D0;
        15'h2940: data = 12'h0D3;
        15'h2941: data = 12'h0D3;
        15'h2942: data = 12'h0D4;
        15'h2943: data = 12'h0D2;
        15'h2944: data = 12'h0D1;
        15'h2945: data = 12'h0CB;
        15'h2946: data = 12'h0C9;
        15'h2947: data = 12'h0C4;
        15'h2948: data = 12'h0C4;
        15'h2949: data = 12'h0BE;
        15'h294A: data = 12'h0B4;
        15'h294B: data = 12'h0B4;
        15'h294C: data = 12'h0AB;
        15'h294D: data = 12'h0AE;
        15'h294E: data = 12'h0AD;
        15'h294F: data = 12'h0AD;
        15'h2950: data = 12'h0B0;
        15'h2951: data = 12'h0B4;
        15'h2952: data = 12'h0AF;
        15'h2953: data = 12'h0A5;
        15'h2954: data = 12'h0A3;
        15'h2955: data = 12'h093;
        15'h2956: data = 12'h086;
        15'h2957: data = 12'h07B;
        15'h2958: data = 12'h071;
        15'h2959: data = 12'h074;
        15'h295A: data = 12'h070;
        15'h295B: data = 12'h072;
        15'h295C: data = 12'h06D;
        15'h295D: data = 12'h06A;
        15'h295E: data = 12'h05F;
        15'h295F: data = 12'h054;
        15'h2960: data = 12'h043;
        15'h2961: data = 12'h7BC;
        15'h2962: data = 12'h7AF;
        15'h2963: data = 12'h7A6;
        15'h2964: data = 12'h7A6;
        15'h2965: data = 12'h79A;
        15'h2966: data = 12'h798;
        15'h2967: data = 12'h78A;
        15'h2968: data = 12'h779;
        15'h2969: data = 12'h76B;
        15'h296A: data = 12'h754;
        15'h296B: data = 12'h743;
        15'h296C: data = 12'h737;
        15'h296D: data = 12'h730;
        15'h296E: data = 12'h729;
        15'h296F: data = 12'h721;
        15'h2970: data = 12'h716;
        15'h2971: data = 12'h70E;
        15'h2972: data = 12'h6FB;
        15'h2973: data = 12'h6E4;
        15'h2974: data = 12'h6D7;
        15'h2975: data = 12'h6C1;
        15'h2976: data = 12'h6B3;
        15'h2977: data = 12'h6A5;
        15'h2978: data = 12'h69A;
        15'h2979: data = 12'h68A;
        15'h297A: data = 12'h681;
        15'h297B: data = 12'h675;
        15'h297C: data = 12'h664;
        15'h297D: data = 12'h659;
        15'h297E: data = 12'h643;
        15'h297F: data = 12'h62F;
        15'h2980: data = 12'h626;
        15'h2981: data = 12'h60A;
        15'h2982: data = 12'h5F5;
        15'h2983: data = 12'h5E4;
        15'h2984: data = 12'h5CB;
        15'h2985: data = 12'h5BD;
        15'h2986: data = 12'h5B1;
        15'h2987: data = 12'h5A3;
        15'h2988: data = 12'h593;
        15'h2989: data = 12'h586;
        15'h298A: data = 12'h574;
        15'h298B: data = 12'h566;
        15'h298C: data = 12'h553;
        15'h298D: data = 12'h543;
        15'h298E: data = 12'h52A;
        15'h298F: data = 12'h518;
        15'h2990: data = 12'h503;
        15'h2991: data = 12'h4F0;
        15'h2992: data = 12'h4D7;
        15'h2993: data = 12'h4C2;
        15'h2994: data = 12'h4AA;
        15'h2995: data = 12'h493;
        15'h2996: data = 12'h47B;
        15'h2997: data = 12'h467;
        15'h2998: data = 12'h44F;
        15'h2999: data = 12'h43F;
        15'h299A: data = 12'h42E;
        15'h299B: data = 12'h417;
        15'h299C: data = 12'h3FF;
        15'h299D: data = 12'h3EC;
        15'h299E: data = 12'h3D9;
        15'h299F: data = 12'h3C3;
        15'h29A0: data = 12'h3B1;
        15'h29A1: data = 12'h397;
        15'h29A2: data = 12'h385;
        15'h29A3: data = 12'h370;
        15'h29A4: data = 12'h35A;
        15'h29A5: data = 12'h346;
        15'h29A6: data = 12'h32F;
        15'h29A7: data = 12'h31C;
        15'h29A8: data = 12'h304;
        15'h29A9: data = 12'h2EF;
        15'h29AA: data = 12'h2DD;
        15'h29AB: data = 12'h2C5;
        15'h29AC: data = 12'h2AA;
        15'h29AD: data = 12'h292;
        15'h29AE: data = 12'h280;
        15'h29AF: data = 12'h266;
        15'h29B0: data = 12'h24F;
        15'h29B1: data = 12'h238;
        15'h29B2: data = 12'h21D;
        15'h29B3: data = 12'h206;
        15'h29B4: data = 12'h1F6;
        15'h29B5: data = 12'h1DA;
        15'h29B6: data = 12'h1C1;
        15'h29B7: data = 12'h1AB;
        15'h29B8: data = 12'h193;
        15'h29B9: data = 12'h17C;
        15'h29BA: data = 12'h166;
        15'h29BB: data = 12'h14E;
        15'h29BC: data = 12'h137;
        15'h29BD: data = 12'h11C;
        15'h29BE: data = 12'h108;
        15'h29BF: data = 12'h0F1;
        15'h29C0: data = 12'h0D9;
        15'h29C1: data = 12'h0BF;
        15'h29C2: data = 12'h0A8;
        15'h29C3: data = 12'h094;
        15'h29C4: data = 12'h080;
        15'h29C5: data = 12'h063;
        15'h29C6: data = 12'h04A;
        15'h29C7: data = 12'h7DF;
        15'h29C8: data = 12'h7CD;
        15'h29C9: data = 12'h7BA;
        15'h29CA: data = 12'h7A3;
        15'h29CB: data = 12'h78B;
        15'h29CC: data = 12'h773;
        15'h29CD: data = 12'h758;
        15'h29CE: data = 12'h748;
        15'h29CF: data = 12'h731;
        15'h29D0: data = 12'h71B;
        15'h29D1: data = 12'h708;
        15'h29D2: data = 12'h6E8;
        15'h29D3: data = 12'h6D7;
        15'h29D4: data = 12'h6BF;
        15'h29D5: data = 12'h6AA;
        15'h29D6: data = 12'h692;
        15'h29D7: data = 12'h67E;
        15'h29D8: data = 12'h662;
        15'h29D9: data = 12'h651;
        15'h29DA: data = 12'h639;
        15'h29DB: data = 12'h627;
        15'h29DC: data = 12'h60D;
        15'h29DD: data = 12'h5F4;
        15'h29DE: data = 12'h5DE;
        15'h29DF: data = 12'h5C7;
        15'h29E0: data = 12'h5B3;
        15'h29E1: data = 12'h59A;
        15'h29E2: data = 12'h582;
        15'h29E3: data = 12'h56D;
        15'h29E4: data = 12'h55D;
        15'h29E5: data = 12'h548;
        15'h29E6: data = 12'h532;
        15'h29E7: data = 12'h519;
        15'h29E8: data = 12'h509;
        15'h29E9: data = 12'h4F3;
        15'h29EA: data = 12'h4E1;
        15'h29EB: data = 12'h4CD;
        15'h29EC: data = 12'h4B8;
        15'h29ED: data = 12'h4A7;
        15'h29EE: data = 12'h497;
        15'h29EF: data = 12'h485;
        15'h29F0: data = 12'h470;
        15'h29F1: data = 12'h45F;
        15'h29F2: data = 12'h44F;
        15'h29F3: data = 12'h445;
        15'h29F4: data = 12'h42F;
        15'h29F5: data = 12'h41E;
        15'h29F6: data = 12'h408;
        15'h29F7: data = 12'h3F9;
        15'h29F8: data = 12'h3E9;
        15'h29F9: data = 12'h3D2;
        15'h29FA: data = 12'h3C0;
        15'h29FB: data = 12'h3AD;
        15'h29FC: data = 12'h398;
        15'h29FD: data = 12'h38C;
        15'h29FE: data = 12'h370;
        15'h29FF: data = 12'h35D;
        15'h2A00: data = 12'h34D;
        15'h2A01: data = 12'h33E;
        15'h2A02: data = 12'h32A;
        15'h2A03: data = 12'h31C;
        15'h2A04: data = 12'h310;
        15'h2A05: data = 12'h300;
        15'h2A06: data = 12'h2F7;
        15'h2A07: data = 12'h2E6;
        15'h2A08: data = 12'h2D8;
        15'h2A09: data = 12'h2D8;
        15'h2A0A: data = 12'h2C9;
        15'h2A0B: data = 12'h2BA;
        15'h2A0C: data = 12'h2AD;
        15'h2A0D: data = 12'h2A1;
        15'h2A0E: data = 12'h294;
        15'h2A0F: data = 12'h280;
        15'h2A10: data = 12'h276;
        15'h2A11: data = 12'h265;
        15'h2A12: data = 12'h259;
        15'h2A13: data = 12'h244;
        15'h2A14: data = 12'h23C;
        15'h2A15: data = 12'h22B;
        15'h2A16: data = 12'h224;
        15'h2A17: data = 12'h216;
        15'h2A18: data = 12'h212;
        15'h2A19: data = 12'h20F;
        15'h2A1A: data = 12'h20F;
        15'h2A1B: data = 12'h1FD;
        15'h2A1C: data = 12'h1FC;
        15'h2A1D: data = 12'h1F2;
        15'h2A1E: data = 12'h1E8;
        15'h2A1F: data = 12'h1E1;
        15'h2A20: data = 12'h1D5;
        15'h2A21: data = 12'h1C7;
        15'h2A22: data = 12'h1BD;
        15'h2A23: data = 12'h1B6;
        15'h2A24: data = 12'h1AA;
        15'h2A25: data = 12'h1A0;
        15'h2A26: data = 12'h197;
        15'h2A27: data = 12'h194;
        15'h2A28: data = 12'h195;
        15'h2A29: data = 12'h193;
        15'h2A2A: data = 12'h191;
        15'h2A2B: data = 12'h190;
        15'h2A2C: data = 12'h18E;
        15'h2A2D: data = 12'h187;
        15'h2A2E: data = 12'h185;
        15'h2A2F: data = 12'h17F;
        15'h2A30: data = 12'h17C;
        15'h2A31: data = 12'h171;
        15'h2A32: data = 12'h16C;
        15'h2A33: data = 12'h169;
        15'h2A34: data = 12'h160;
        15'h2A35: data = 12'h15D;
        15'h2A36: data = 12'h160;
        15'h2A37: data = 12'h162;
        15'h2A38: data = 12'h15C;
        15'h2A39: data = 12'h160;
        15'h2A3A: data = 12'h163;
        15'h2A3B: data = 12'h16A;
        15'h2A3C: data = 12'h167;
        15'h2A3D: data = 12'h169;
        15'h2A3E: data = 12'h169;
        15'h2A3F: data = 12'h16E;
        15'h2A40: data = 12'h16C;
        15'h2A41: data = 12'h169;
        15'h2A42: data = 12'h162;
        15'h2A43: data = 12'h15E;
        15'h2A44: data = 12'h166;
        15'h2A45: data = 12'h164;
        15'h2A46: data = 12'h16A;
        15'h2A47: data = 12'h16C;
        15'h2A48: data = 12'h16F;
        15'h2A49: data = 12'h17E;
        15'h2A4A: data = 12'h188;
        15'h2A4B: data = 12'h18D;
        15'h2A4C: data = 12'h195;
        15'h2A4D: data = 12'h197;
        15'h2A4E: data = 12'h19E;
        15'h2A4F: data = 12'h1A4;
        15'h2A50: data = 12'h1A8;
        15'h2A51: data = 12'h1B0;
        15'h2A52: data = 12'h1B1;
        15'h2A53: data = 12'h1AF;
        15'h2A54: data = 12'h1B6;
        15'h2A55: data = 12'h1BE;
        15'h2A56: data = 12'h1C1;
        15'h2A57: data = 12'h1CC;
        15'h2A58: data = 12'h1D1;
        15'h2A59: data = 12'h1D8;
        15'h2A5A: data = 12'h1E9;
        15'h2A5B: data = 12'h1FB;
        15'h2A5C: data = 12'h205;
        15'h2A5D: data = 12'h211;
        15'h2A5E: data = 12'h220;
        15'h2A5F: data = 12'h224;
        15'h2A60: data = 12'h232;
        15'h2A61: data = 12'h237;
        15'h2A62: data = 12'h245;
        15'h2A63: data = 12'h247;
        15'h2A64: data = 12'h255;
        15'h2A65: data = 12'h258;
        15'h2A66: data = 12'h264;
        15'h2A67: data = 12'h26E;
        15'h2A68: data = 12'h27B;
        15'h2A69: data = 12'h288;
        15'h2A6A: data = 12'h294;
        15'h2A6B: data = 12'h2A6;
        15'h2A6C: data = 12'h2B7;
        15'h2A6D: data = 12'h2C9;
        15'h2A6E: data = 12'h2DF;
        15'h2A6F: data = 12'h2E9;
        15'h2A70: data = 12'h2FA;
        15'h2A71: data = 12'h309;
        15'h2A72: data = 12'h31A;
        15'h2A73: data = 12'h329;
        15'h2A74: data = 12'h338;
        15'h2A75: data = 12'h345;
        15'h2A76: data = 12'h351;
        15'h2A77: data = 12'h35E;
        15'h2A78: data = 12'h36A;
        15'h2A79: data = 12'h373;
        15'h2A7A: data = 12'h38D;
        15'h2A7B: data = 12'h391;
        15'h2A7C: data = 12'h3A4;
        15'h2A7D: data = 12'h3B7;
        15'h2A7E: data = 12'h3C9;
        15'h2A7F: data = 12'h3DD;
        15'h2A80: data = 12'h3F1;
        15'h2A81: data = 12'h404;
        15'h2A82: data = 12'h421;
        15'h2A83: data = 12'h432;
        15'h2A84: data = 12'h44B;
        15'h2A85: data = 12'h45E;
        15'h2A86: data = 12'h46C;
        15'h2A87: data = 12'h485;
        15'h2A88: data = 12'h493;
        15'h2A89: data = 12'h4A8;
        15'h2A8A: data = 12'h4B8;
        15'h2A8B: data = 12'h4CD;
        15'h2A8C: data = 12'h4DF;
        15'h2A8D: data = 12'h4ED;
        15'h2A8E: data = 12'h4FF;
        15'h2A8F: data = 12'h513;
        15'h2A90: data = 12'h523;
        15'h2A91: data = 12'h53C;
        15'h2A92: data = 12'h551;
        15'h2A93: data = 12'h568;
        15'h2A94: data = 12'h579;
        15'h2A95: data = 12'h58D;
        15'h2A96: data = 12'h5A6;
        15'h2A97: data = 12'h5BC;
        15'h2A98: data = 12'h5D4;
        15'h2A99: data = 12'h5EC;
        15'h2A9A: data = 12'h608;
        15'h2A9B: data = 12'h621;
        15'h2A9C: data = 12'h636;
        15'h2A9D: data = 12'h64B;
        15'h2A9E: data = 12'h664;
        15'h2A9F: data = 12'h679;
        15'h2AA0: data = 12'h691;
        15'h2AA1: data = 12'h69F;
        15'h2AA2: data = 12'h6B5;
        15'h2AA3: data = 12'h6C9;
        15'h2AA4: data = 12'h6DE;
        15'h2AA5: data = 12'h6F0;
        15'h2AA6: data = 12'h707;
        15'h2AA7: data = 12'h718;
        15'h2AA8: data = 12'h733;
        15'h2AA9: data = 12'h743;
        15'h2AAA: data = 12'h75A;
        15'h2AAB: data = 12'h775;
        15'h2AAC: data = 12'h792;
        15'h2AAD: data = 12'h7A3;
        15'h2AAE: data = 12'h7C0;
        15'h2AAF: data = 12'h7DB;
        15'h2AB0: data = 12'h7F3;
        15'h2AB1: data = 12'h806;
        15'h2AB2: data = 12'h079;
        15'h2AB3: data = 12'h090;
        15'h2AB4: data = 12'h0A5;
        15'h2AB5: data = 12'h0B9;
        15'h2AB6: data = 12'h0D6;
        15'h2AB7: data = 12'h0EC;
        15'h2AB8: data = 12'h0FE;
        15'h2AB9: data = 12'h111;
        15'h2ABA: data = 12'h128;
        15'h2ABB: data = 12'h140;
        15'h2ABC: data = 12'h152;
        15'h2ABD: data = 12'h167;
        15'h2ABE: data = 12'h178;
        15'h2ABF: data = 12'h192;
        15'h2AC0: data = 12'h1A9;
        15'h2AC1: data = 12'h1BB;
        15'h2AC2: data = 12'h1D3;
        15'h2AC3: data = 12'h1EB;
        15'h2AC4: data = 12'h204;
        15'h2AC5: data = 12'h219;
        15'h2AC6: data = 12'h232;
        15'h2AC7: data = 12'h24C;
        15'h2AC8: data = 12'h262;
        15'h2AC9: data = 12'h279;
        15'h2ACA: data = 12'h295;
        15'h2ACB: data = 12'h2AE;
        15'h2ACC: data = 12'h2C6;
        15'h2ACD: data = 12'h2DB;
        15'h2ACE: data = 12'h2F5;
        15'h2ACF: data = 12'h30B;
        15'h2AD0: data = 12'h327;
        15'h2AD1: data = 12'h33B;
        15'h2AD2: data = 12'h350;
        15'h2AD3: data = 12'h36C;
        15'h2AD4: data = 12'h37E;
        15'h2AD5: data = 12'h39B;
        15'h2AD6: data = 12'h3AA;
        15'h2AD7: data = 12'h3C3;
        15'h2AD8: data = 12'h3D7;
        15'h2AD9: data = 12'h3EE;
        15'h2ADA: data = 12'h3FF;
        15'h2ADB: data = 12'h415;
        15'h2ADC: data = 12'h429;
        15'h2ADD: data = 12'h441;
        15'h2ADE: data = 12'h44B;
        15'h2ADF: data = 12'h462;
        15'h2AE0: data = 12'h476;
        15'h2AE1: data = 12'h48F;
        15'h2AE2: data = 12'h4A1;
        15'h2AE3: data = 12'h4B0;
        15'h2AE4: data = 12'h4C0;
        15'h2AE5: data = 12'h4D5;
        15'h2AE6: data = 12'h4ED;
        15'h2AE7: data = 12'h503;
        15'h2AE8: data = 12'h50D;
        15'h2AE9: data = 12'h523;
        15'h2AEA: data = 12'h538;
        15'h2AEB: data = 12'h547;
        15'h2AEC: data = 12'h55B;
        15'h2AED: data = 12'h56B;
        15'h2AEE: data = 12'h584;
        15'h2AEF: data = 12'h592;
        15'h2AF0: data = 12'h5A9;
        15'h2AF1: data = 12'h5BA;
        15'h2AF2: data = 12'h5C7;
        15'h2AF3: data = 12'h5DA;
        15'h2AF4: data = 12'h5F1;
        15'h2AF5: data = 12'h603;
        15'h2AF6: data = 12'h610;
        15'h2AF7: data = 12'h620;
        15'h2AF8: data = 12'h634;
        15'h2AF9: data = 12'h642;
        15'h2AFA: data = 12'h658;
        15'h2AFB: data = 12'h668;
        15'h2AFC: data = 12'h679;
        15'h2AFD: data = 12'h687;
        15'h2AFE: data = 12'h69B;
        15'h2AFF: data = 12'h6A8;
        15'h2B00: data = 12'h6B8;
        15'h2B01: data = 12'h6C9;
        15'h2B02: data = 12'h6D8;
        15'h2B03: data = 12'h6DE;
        15'h2B04: data = 12'h6EF;
        15'h2B05: data = 12'h6FF;
        15'h2B06: data = 12'h709;
        15'h2B07: data = 12'h717;
        15'h2B08: data = 12'h723;
        15'h2B09: data = 12'h737;
        15'h2B0A: data = 12'h73A;
        15'h2B0B: data = 12'h744;
        15'h2B0C: data = 12'h753;
        15'h2B0D: data = 12'h75D;
        15'h2B0E: data = 12'h766;
        15'h2B0F: data = 12'h776;
        15'h2B10: data = 12'h77F;
        15'h2B11: data = 12'h78D;
        15'h2B12: data = 12'h793;
        15'h2B13: data = 12'h79B;
        15'h2B14: data = 12'h7A1;
        15'h2B15: data = 12'h7AC;
        15'h2B16: data = 12'h7B4;
        15'h2B17: data = 12'h7BD;
        15'h2B18: data = 12'h7C1;
        15'h2B19: data = 12'h7C5;
        15'h2B1A: data = 12'h7CD;
        15'h2B1B: data = 12'h7D4;
        15'h2B1C: data = 12'h7E1;
        15'h2B1D: data = 12'h7E6;
        15'h2B1E: data = 12'h7EC;
        15'h2B1F: data = 12'h7EF;
        15'h2B20: data = 12'h7F8;
        15'h2B21: data = 12'h7FA;
        15'h2B22: data = 12'h7FD;
        15'h2B23: data = 12'h805;
        15'h2B24: data = 12'h62C;
        15'h2B25: data = 12'h083;
        15'h2B26: data = 12'h092;
        15'h2B27: data = 12'h094;
        15'h2B28: data = 12'h096;
        15'h2B29: data = 12'h09E;
        15'h2B2A: data = 12'h09F;
        15'h2B2B: data = 12'h0AB;
        15'h2B2C: data = 12'h0AA;
        15'h2B2D: data = 12'h0AD;
        15'h2B2E: data = 12'h0B8;
        15'h2B2F: data = 12'h0B9;
        15'h2B30: data = 12'h0BB;
        15'h2B31: data = 12'h0BC;
        15'h2B32: data = 12'h0CB;
        15'h2B33: data = 12'h0D0;
        15'h2B34: data = 12'h0CF;
        15'h2B35: data = 12'h0D2;
        15'h2B36: data = 12'h0D7;
        15'h2B37: data = 12'h0D3;
        15'h2B38: data = 12'h0D7;
        15'h2B39: data = 12'h0CB;
        15'h2B3A: data = 12'h0CB;
        15'h2B3B: data = 12'h0C8;
        15'h2B3C: data = 12'h0C6;
        15'h2B3D: data = 12'h0BF;
        15'h2B3E: data = 12'h0B4;
        15'h2B3F: data = 12'h0B6;
        15'h2B40: data = 12'h0AD;
        15'h2B41: data = 12'h0AE;
        15'h2B42: data = 12'h0A8;
        15'h2B43: data = 12'h0AC;
        15'h2B44: data = 12'h0B0;
        15'h2B45: data = 12'h0B3;
        15'h2B46: data = 12'h0AB;
        15'h2B47: data = 12'h0A3;
        15'h2B48: data = 12'h0A4;
        15'h2B49: data = 12'h097;
        15'h2B4A: data = 12'h08A;
        15'h2B4B: data = 12'h07D;
        15'h2B4C: data = 12'h075;
        15'h2B4D: data = 12'h075;
        15'h2B4E: data = 12'h072;
        15'h2B4F: data = 12'h06F;
        15'h2B50: data = 12'h06B;
        15'h2B51: data = 12'h067;
        15'h2B52: data = 12'h05E;
        15'h2B53: data = 12'h055;
        15'h2B54: data = 12'h043;
        15'h2B55: data = 12'h7BB;
        15'h2B56: data = 12'h7AF;
        15'h2B57: data = 12'h7A8;
        15'h2B58: data = 12'h7A1;
        15'h2B59: data = 12'h79C;
        15'h2B5A: data = 12'h793;
        15'h2B5B: data = 12'h789;
        15'h2B5C: data = 12'h776;
        15'h2B5D: data = 12'h76A;
        15'h2B5E: data = 12'h751;
        15'h2B5F: data = 12'h744;
        15'h2B60: data = 12'h735;
        15'h2B61: data = 12'h72E;
        15'h2B62: data = 12'h725;
        15'h2B63: data = 12'h71D;
        15'h2B64: data = 12'h715;
        15'h2B65: data = 12'h705;
        15'h2B66: data = 12'h6FA;
        15'h2B67: data = 12'h6E6;
        15'h2B68: data = 12'h6D8;
        15'h2B69: data = 12'h6C7;
        15'h2B6A: data = 12'h6B2;
        15'h2B6B: data = 12'h6A6;
        15'h2B6C: data = 12'h696;
        15'h2B6D: data = 12'h688;
        15'h2B6E: data = 12'h67D;
        15'h2B6F: data = 12'h672;
        15'h2B70: data = 12'h667;
        15'h2B71: data = 12'h657;
        15'h2B72: data = 12'h646;
        15'h2B73: data = 12'h632;
        15'h2B74: data = 12'h628;
        15'h2B75: data = 12'h60A;
        15'h2B76: data = 12'h5F7;
        15'h2B77: data = 12'h5E5;
        15'h2B78: data = 12'h5CA;
        15'h2B79: data = 12'h5BD;
        15'h2B7A: data = 12'h5B0;
        15'h2B7B: data = 12'h5A0;
        15'h2B7C: data = 12'h58F;
        15'h2B7D: data = 12'h581;
        15'h2B7E: data = 12'h572;
        15'h2B7F: data = 12'h564;
        15'h2B80: data = 12'h556;
        15'h2B81: data = 12'h542;
        15'h2B82: data = 12'h52F;
        15'h2B83: data = 12'h519;
        15'h2B84: data = 12'h505;
        15'h2B85: data = 12'h4F2;
        15'h2B86: data = 12'h4D5;
        15'h2B87: data = 12'h4C0;
        15'h2B88: data = 12'h4AD;
        15'h2B89: data = 12'h495;
        15'h2B8A: data = 12'h47E;
        15'h2B8B: data = 12'h46B;
        15'h2B8C: data = 12'h452;
        15'h2B8D: data = 12'h43D;
        15'h2B8E: data = 12'h429;
        15'h2B8F: data = 12'h416;
        15'h2B90: data = 12'h401;
        15'h2B91: data = 12'h3EA;
        15'h2B92: data = 12'h3D4;
        15'h2B93: data = 12'h3C1;
        15'h2B94: data = 12'h3B1;
        15'h2B95: data = 12'h392;
        15'h2B96: data = 12'h383;
        15'h2B97: data = 12'h369;
        15'h2B98: data = 12'h356;
        15'h2B99: data = 12'h341;
        15'h2B9A: data = 12'h331;
        15'h2B9B: data = 12'h31D;
        15'h2B9C: data = 12'h303;
        15'h2B9D: data = 12'h2EE;
        15'h2B9E: data = 12'h2D9;
        15'h2B9F: data = 12'h2C3;
        15'h2BA0: data = 12'h2AB;
        15'h2BA1: data = 12'h290;
        15'h2BA2: data = 12'h27F;
        15'h2BA3: data = 12'h265;
        15'h2BA4: data = 12'h249;
        15'h2BA5: data = 12'h238;
        15'h2BA6: data = 12'h21E;
        15'h2BA7: data = 12'h205;
        15'h2BA8: data = 12'h1F4;
        15'h2BA9: data = 12'h1D9;
        15'h2BAA: data = 12'h1C2;
        15'h2BAB: data = 12'h1A9;
        15'h2BAC: data = 12'h193;
        15'h2BAD: data = 12'h17D;
        15'h2BAE: data = 12'h164;
        15'h2BAF: data = 12'h14D;
        15'h2BB0: data = 12'h135;
        15'h2BB1: data = 12'h11E;
        15'h2BB2: data = 12'h10A;
        15'h2BB3: data = 12'h0F3;
        15'h2BB4: data = 12'h0DB;
        15'h2BB5: data = 12'h0C1;
        15'h2BB6: data = 12'h0A4;
        15'h2BB7: data = 12'h08D;
        15'h2BB8: data = 12'h07C;
        15'h2BB9: data = 12'h063;
        15'h2BBA: data = 12'h04A;
        15'h2BBB: data = 12'h7DD;
        15'h2BBC: data = 12'h7CC;
        15'h2BBD: data = 12'h7B5;
        15'h2BBE: data = 12'h7A2;
        15'h2BBF: data = 12'h789;
        15'h2BC0: data = 12'h774;
        15'h2BC1: data = 12'h759;
        15'h2BC2: data = 12'h745;
        15'h2BC3: data = 12'h733;
        15'h2BC4: data = 12'h71C;
        15'h2BC5: data = 12'h705;
        15'h2BC6: data = 12'h6EA;
        15'h2BC7: data = 12'h6D4;
        15'h2BC8: data = 12'h6C1;
        15'h2BC9: data = 12'h6A8;
        15'h2BCA: data = 12'h693;
        15'h2BCB: data = 12'h67E;
        15'h2BCC: data = 12'h665;
        15'h2BCD: data = 12'h651;
        15'h2BCE: data = 12'h636;
        15'h2BCF: data = 12'h627;
        15'h2BD0: data = 12'h60F;
        15'h2BD1: data = 12'h5F6;
        15'h2BD2: data = 12'h5E0;
        15'h2BD3: data = 12'h5C7;
        15'h2BD4: data = 12'h5B5;
        15'h2BD5: data = 12'h597;
        15'h2BD6: data = 12'h582;
        15'h2BD7: data = 12'h56B;
        15'h2BD8: data = 12'h558;
        15'h2BD9: data = 12'h545;
        15'h2BDA: data = 12'h532;
        15'h2BDB: data = 12'h51D;
        15'h2BDC: data = 12'h507;
        15'h2BDD: data = 12'h4F4;
        15'h2BDE: data = 12'h4DC;
        15'h2BDF: data = 12'h4CD;
        15'h2BE0: data = 12'h4B6;
        15'h2BE1: data = 12'h4A3;
        15'h2BE2: data = 12'h492;
        15'h2BE3: data = 12'h480;
        15'h2BE4: data = 12'h46F;
        15'h2BE5: data = 12'h45D;
        15'h2BE6: data = 12'h450;
        15'h2BE7: data = 12'h43F;
        15'h2BE8: data = 12'h42C;
        15'h2BE9: data = 12'h419;
        15'h2BEA: data = 12'h407;
        15'h2BEB: data = 12'h3FC;
        15'h2BEC: data = 12'h3EB;
        15'h2BED: data = 12'h3D3;
        15'h2BEE: data = 12'h3C0;
        15'h2BEF: data = 12'h3AC;
        15'h2BF0: data = 12'h39A;
        15'h2BF1: data = 12'h390;
        15'h2BF2: data = 12'h375;
        15'h2BF3: data = 12'h361;
        15'h2BF4: data = 12'h34E;
        15'h2BF5: data = 12'h33D;
        15'h2BF6: data = 12'h32E;
        15'h2BF7: data = 12'h31C;
        15'h2BF8: data = 12'h30E;
        15'h2BF9: data = 12'h2FE;
        15'h2BFA: data = 12'h2F2;
        15'h2BFB: data = 12'h2E4;
        15'h2BFC: data = 12'h2DC;
        15'h2BFD: data = 12'h2D7;
        15'h2BFE: data = 12'h2CA;
        15'h2BFF: data = 12'h2BB;
        15'h2C00: data = 12'h2AE;
        15'h2C01: data = 12'h2A1;
        15'h2C02: data = 12'h294;
        15'h2C03: data = 12'h283;
        15'h2C04: data = 12'h27C;
        15'h2C05: data = 12'h262;
        15'h2C06: data = 12'h25A;
        15'h2C07: data = 12'h248;
        15'h2C08: data = 12'h240;
        15'h2C09: data = 12'h22D;
        15'h2C0A: data = 12'h225;
        15'h2C0B: data = 12'h21B;
        15'h2C0C: data = 12'h214;
        15'h2C0D: data = 12'h20E;
        15'h2C0E: data = 12'h209;
        15'h2C0F: data = 12'h1FD;
        15'h2C10: data = 12'h1F7;
        15'h2C11: data = 12'h1EF;
        15'h2C12: data = 12'h1EB;
        15'h2C13: data = 12'h1DE;
        15'h2C14: data = 12'h1D2;
        15'h2C15: data = 12'h1C7;
        15'h2C16: data = 12'h1BB;
        15'h2C17: data = 12'h1B3;
        15'h2C18: data = 12'h1A9;
        15'h2C19: data = 12'h1A0;
        15'h2C1A: data = 12'h19A;
        15'h2C1B: data = 12'h194;
        15'h2C1C: data = 12'h193;
        15'h2C1D: data = 12'h191;
        15'h2C1E: data = 12'h18C;
        15'h2C1F: data = 12'h18F;
        15'h2C20: data = 12'h18E;
        15'h2C21: data = 12'h186;
        15'h2C22: data = 12'h187;
        15'h2C23: data = 12'h17C;
        15'h2C24: data = 12'h17B;
        15'h2C25: data = 12'h172;
        15'h2C26: data = 12'h170;
        15'h2C27: data = 12'h169;
        15'h2C28: data = 12'h160;
        15'h2C29: data = 12'h15D;
        15'h2C2A: data = 12'h15D;
        15'h2C2B: data = 12'h15E;
        15'h2C2C: data = 12'h159;
        15'h2C2D: data = 12'h15C;
        15'h2C2E: data = 12'h15F;
        15'h2C2F: data = 12'h165;
        15'h2C30: data = 12'h165;
        15'h2C31: data = 12'h168;
        15'h2C32: data = 12'h169;
        15'h2C33: data = 12'h16D;
        15'h2C34: data = 12'h16E;
        15'h2C35: data = 12'h169;
        15'h2C36: data = 12'h165;
        15'h2C37: data = 12'h164;
        15'h2C38: data = 12'h167;
        15'h2C39: data = 12'h164;
        15'h2C3A: data = 12'h168;
        15'h2C3B: data = 12'h16D;
        15'h2C3C: data = 12'h16E;
        15'h2C3D: data = 12'h17B;
        15'h2C3E: data = 12'h187;
        15'h2C3F: data = 12'h18B;
        15'h2C40: data = 12'h195;
        15'h2C41: data = 12'h193;
        15'h2C42: data = 12'h19F;
        15'h2C43: data = 12'h1A4;
        15'h2C44: data = 12'h1AD;
        15'h2C45: data = 12'h1B1;
        15'h2C46: data = 12'h1AD;
        15'h2C47: data = 12'h1AF;
        15'h2C48: data = 12'h1B7;
        15'h2C49: data = 12'h1BA;
        15'h2C4A: data = 12'h1C1;
        15'h2C4B: data = 12'h1C9;
        15'h2C4C: data = 12'h1D2;
        15'h2C4D: data = 12'h1DA;
        15'h2C4E: data = 12'h1E6;
        15'h2C4F: data = 12'h1FA;
        15'h2C50: data = 12'h204;
        15'h2C51: data = 12'h210;
        15'h2C52: data = 12'h21F;
        15'h2C53: data = 12'h221;
        15'h2C54: data = 12'h22E;
        15'h2C55: data = 12'h238;
        15'h2C56: data = 12'h247;
        15'h2C57: data = 12'h24C;
        15'h2C58: data = 12'h258;
        15'h2C59: data = 12'h25A;
        15'h2C5A: data = 12'h268;
        15'h2C5B: data = 12'h269;
        15'h2C5C: data = 12'h27A;
        15'h2C5D: data = 12'h286;
        15'h2C5E: data = 12'h294;
        15'h2C5F: data = 12'h2A2;
        15'h2C60: data = 12'h2B6;
        15'h2C61: data = 12'h2C5;
        15'h2C62: data = 12'h2D8;
        15'h2C63: data = 12'h2E6;
        15'h2C64: data = 12'h2F8;
        15'h2C65: data = 12'h308;
        15'h2C66: data = 12'h31B;
        15'h2C67: data = 12'h327;
        15'h2C68: data = 12'h335;
        15'h2C69: data = 12'h345;
        15'h2C6A: data = 12'h357;
        15'h2C6B: data = 12'h361;
        15'h2C6C: data = 12'h36D;
        15'h2C6D: data = 12'h378;
        15'h2C6E: data = 12'h38D;
        15'h2C6F: data = 12'h393;
        15'h2C70: data = 12'h3A7;
        15'h2C71: data = 12'h3B6;
        15'h2C72: data = 12'h3C7;
        15'h2C73: data = 12'h3DD;
        15'h2C74: data = 12'h3F1;
        15'h2C75: data = 12'h401;
        15'h2C76: data = 12'h41C;
        15'h2C77: data = 12'h431;
        15'h2C78: data = 12'h447;
        15'h2C79: data = 12'h45A;
        15'h2C7A: data = 12'h46D;
        15'h2C7B: data = 12'h482;
        15'h2C7C: data = 12'h493;
        15'h2C7D: data = 12'h4AB;
        15'h2C7E: data = 12'h4BA;
        15'h2C7F: data = 12'h4CE;
        15'h2C80: data = 12'h4E1;
        15'h2C81: data = 12'h4F3;
        15'h2C82: data = 12'h508;
        15'h2C83: data = 12'h516;
        15'h2C84: data = 12'h525;
        15'h2C85: data = 12'h53A;
        15'h2C86: data = 12'h550;
        15'h2C87: data = 12'h565;
        15'h2C88: data = 12'h573;
        15'h2C89: data = 12'h58C;
        15'h2C8A: data = 12'h5A4;
        15'h2C8B: data = 12'h5BB;
        15'h2C8C: data = 12'h5D2;
        15'h2C8D: data = 12'h5EF;
        15'h2C8E: data = 12'h605;
        15'h2C8F: data = 12'h61D;
        15'h2C90: data = 12'h637;
        15'h2C91: data = 12'h64B;
        15'h2C92: data = 12'h663;
        15'h2C93: data = 12'h678;
        15'h2C94: data = 12'h691;
        15'h2C95: data = 12'h6A1;
        15'h2C96: data = 12'h6B5;
        15'h2C97: data = 12'h6CB;
        15'h2C98: data = 12'h6DC;
        15'h2C99: data = 12'h6F0;
        15'h2C9A: data = 12'h703;
        15'h2C9B: data = 12'h716;
        15'h2C9C: data = 12'h732;
        15'h2C9D: data = 12'h744;
        15'h2C9E: data = 12'h756;
        15'h2C9F: data = 12'h772;
        15'h2CA0: data = 12'h78F;
        15'h2CA1: data = 12'h7A2;
        15'h2CA2: data = 12'h7BD;
        15'h2CA3: data = 12'h7D9;
        15'h2CA4: data = 12'h7F0;
        15'h2CA5: data = 12'h80A;
        15'h2CA6: data = 12'h0A5;
        15'h2CA7: data = 12'h090;
        15'h2CA8: data = 12'h0A5;
        15'h2CA9: data = 12'h0BA;
        15'h2CAA: data = 12'h0D2;
        15'h2CAB: data = 12'h0E9;
        15'h2CAC: data = 12'h101;
        15'h2CAD: data = 12'h115;
        15'h2CAE: data = 12'h12B;
        15'h2CAF: data = 12'h140;
        15'h2CB0: data = 12'h151;
        15'h2CB1: data = 12'h167;
        15'h2CB2: data = 12'h17C;
        15'h2CB3: data = 12'h196;
        15'h2CB4: data = 12'h1AD;
        15'h2CB5: data = 12'h1BD;
        15'h2CB6: data = 12'h1D4;
        15'h2CB7: data = 12'h1EF;
        15'h2CB8: data = 12'h206;
        15'h2CB9: data = 12'h216;
        15'h2CBA: data = 12'h233;
        15'h2CBB: data = 12'h24B;
        15'h2CBC: data = 12'h266;
        15'h2CBD: data = 12'h279;
        15'h2CBE: data = 12'h28F;
        15'h2CBF: data = 12'h2AA;
        15'h2CC0: data = 12'h2C7;
        15'h2CC1: data = 12'h2DE;
        15'h2CC2: data = 12'h2F7;
        15'h2CC3: data = 12'h30F;
        15'h2CC4: data = 12'h329;
        15'h2CC5: data = 12'h33A;
        15'h2CC6: data = 12'h34F;
        15'h2CC7: data = 12'h369;
        15'h2CC8: data = 12'h380;
        15'h2CC9: data = 12'h39C;
        15'h2CCA: data = 12'h3AC;
        15'h2CCB: data = 12'h3C0;
        15'h2CCC: data = 12'h3D9;
        15'h2CCD: data = 12'h3F1;
        15'h2CCE: data = 12'h3FE;
        15'h2CCF: data = 12'h418;
        15'h2CD0: data = 12'h42D;
        15'h2CD1: data = 12'h442;
        15'h2CD2: data = 12'h453;
        15'h2CD3: data = 12'h467;
        15'h2CD4: data = 12'h47B;
        15'h2CD5: data = 12'h492;
        15'h2CD6: data = 12'h4A6;
        15'h2CD7: data = 12'h4B5;
        15'h2CD8: data = 12'h4C3;
        15'h2CD9: data = 12'h4DA;
        15'h2CDA: data = 12'h4EF;
        15'h2CDB: data = 12'h504;
        15'h2CDC: data = 12'h510;
        15'h2CDD: data = 12'h526;
        15'h2CDE: data = 12'h53A;
        15'h2CDF: data = 12'h547;
        15'h2CE0: data = 12'h55C;
        15'h2CE1: data = 12'h56A;
        15'h2CE2: data = 12'h581;
        15'h2CE3: data = 12'h593;
        15'h2CE4: data = 12'h5A8;
        15'h2CE5: data = 12'h5BB;
        15'h2CE6: data = 12'h5C7;
        15'h2CE7: data = 12'h5D8;
        15'h2CE8: data = 12'h5EE;
        15'h2CE9: data = 12'h601;
        15'h2CEA: data = 12'h60D;
        15'h2CEB: data = 12'h61F;
        15'h2CEC: data = 12'h632;
        15'h2CED: data = 12'h643;
        15'h2CEE: data = 12'h654;
        15'h2CEF: data = 12'h66A;
        15'h2CF0: data = 12'h677;
        15'h2CF1: data = 12'h68A;
        15'h2CF2: data = 12'h69A;
        15'h2CF3: data = 12'h6A9;
        15'h2CF4: data = 12'h6B7;
        15'h2CF5: data = 12'h6C5;
        15'h2CF6: data = 12'h6D8;
        15'h2CF7: data = 12'h6E1;
        15'h2CF8: data = 12'h6EE;
        15'h2CF9: data = 12'h701;
        15'h2CFA: data = 12'h70C;
        15'h2CFB: data = 12'h714;
        15'h2CFC: data = 12'h725;
        15'h2CFD: data = 12'h737;
        15'h2CFE: data = 12'h739;
        15'h2CFF: data = 12'h745;
        15'h2D00: data = 12'h74E;
        15'h2D01: data = 12'h75E;
        15'h2D02: data = 12'h766;
        15'h2D03: data = 12'h775;
        15'h2D04: data = 12'h77D;
        15'h2D05: data = 12'h78B;
        15'h2D06: data = 12'h790;
        15'h2D07: data = 12'h79A;
        15'h2D08: data = 12'h7A2;
        15'h2D09: data = 12'h7AF;
        15'h2D0A: data = 12'h7B6;
        15'h2D0B: data = 12'h7BF;
        15'h2D0C: data = 12'h7C4;
        15'h2D0D: data = 12'h7CB;
        15'h2D0E: data = 12'h7D4;
        15'h2D0F: data = 12'h7D8;
        15'h2D10: data = 12'h7E4;
        15'h2D11: data = 12'h7E5;
        15'h2D12: data = 12'h7EC;
        15'h2D13: data = 12'h7F5;
        15'h2D14: data = 12'h7FB;
        15'h2D15: data = 12'h7FE;
        15'h2D16: data = 12'h7FE;
        15'h2D17: data = 12'h805;
        15'h2D18: data = 12'h634;
        15'h2D19: data = 12'h087;
        15'h2D1A: data = 12'h091;
        15'h2D1B: data = 12'h095;
        15'h2D1C: data = 12'h096;
        15'h2D1D: data = 12'h0A1;
        15'h2D1E: data = 12'h0A3;
        15'h2D1F: data = 12'h0A9;
        15'h2D20: data = 12'h0AE;
        15'h2D21: data = 12'h0AE;
        15'h2D22: data = 12'h0B9;
        15'h2D23: data = 12'h0BC;
        15'h2D24: data = 12'h0BD;
        15'h2D25: data = 12'h0C0;
        15'h2D26: data = 12'h0CB;
        15'h2D27: data = 12'h0CE;
        15'h2D28: data = 12'h0D1;
        15'h2D29: data = 12'h0D5;
        15'h2D2A: data = 12'h0D7;
        15'h2D2B: data = 12'h0D4;
        15'h2D2C: data = 12'h0D5;
        15'h2D2D: data = 12'h0CF;
        15'h2D2E: data = 12'h0CD;
        15'h2D2F: data = 12'h0CB;
        15'h2D30: data = 12'h0C8;
        15'h2D31: data = 12'h0C2;
        15'h2D32: data = 12'h0B9;
        15'h2D33: data = 12'h0B6;
        15'h2D34: data = 12'h0AF;
        15'h2D35: data = 12'h0AF;
        15'h2D36: data = 12'h0A8;
        15'h2D37: data = 12'h0AE;
        15'h2D38: data = 12'h0AD;
        15'h2D39: data = 12'h0B2;
        15'h2D3A: data = 12'h0B0;
        15'h2D3B: data = 12'h0A5;
        15'h2D3C: data = 12'h0A2;
        15'h2D3D: data = 12'h09E;
        15'h2D3E: data = 12'h08E;
        15'h2D3F: data = 12'h081;
        15'h2D40: data = 12'h073;
        15'h2D41: data = 12'h072;
        15'h2D42: data = 12'h070;
        15'h2D43: data = 12'h06E;
        15'h2D44: data = 12'h069;
        15'h2D45: data = 12'h067;
        15'h2D46: data = 12'h05F;
        15'h2D47: data = 12'h053;
        15'h2D48: data = 12'h046;
        15'h2D49: data = 12'h7C0;
        15'h2D4A: data = 12'h7B2;
        15'h2D4B: data = 12'h7A6;
        15'h2D4C: data = 12'h7A0;
        15'h2D4D: data = 12'h79C;
        15'h2D4E: data = 12'h794;
        15'h2D4F: data = 12'h78C;
        15'h2D50: data = 12'h779;
        15'h2D51: data = 12'h76F;
        15'h2D52: data = 12'h75A;
        15'h2D53: data = 12'h743;
        15'h2D54: data = 12'h734;
        15'h2D55: data = 12'h72E;
        15'h2D56: data = 12'h727;
        15'h2D57: data = 12'h71E;
        15'h2D58: data = 12'h712;
        15'h2D59: data = 12'h70F;
        15'h2D5A: data = 12'h6FE;
        15'h2D5B: data = 12'h6EA;
        15'h2D5C: data = 12'h6DC;
        15'h2D5D: data = 12'h6C8;
        15'h2D5E: data = 12'h6B1;
        15'h2D5F: data = 12'h6A3;
        15'h2D60: data = 12'h694;
        15'h2D61: data = 12'h687;
        15'h2D62: data = 12'h67E;
        15'h2D63: data = 12'h676;
        15'h2D64: data = 12'h667;
        15'h2D65: data = 12'h658;
        15'h2D66: data = 12'h646;
        15'h2D67: data = 12'h634;
        15'h2D68: data = 12'h629;
        15'h2D69: data = 12'h60E;
        15'h2D6A: data = 12'h5F9;
        15'h2D6B: data = 12'h5E4;
        15'h2D6C: data = 12'h5CF;
        15'h2D6D: data = 12'h5BF;
        15'h2D6E: data = 12'h5B1;
        15'h2D6F: data = 12'h5A2;
        15'h2D70: data = 12'h592;
        15'h2D71: data = 12'h580;
        15'h2D72: data = 12'h573;
        15'h2D73: data = 12'h564;
        15'h2D74: data = 12'h552;
        15'h2D75: data = 12'h541;
        15'h2D76: data = 12'h52C;
        15'h2D77: data = 12'h519;
        15'h2D78: data = 12'h506;
        15'h2D79: data = 12'h4F3;
        15'h2D7A: data = 12'h4DC;
        15'h2D7B: data = 12'h4C6;
        15'h2D7C: data = 12'h4B1;
        15'h2D7D: data = 12'h496;
        15'h2D7E: data = 12'h47E;
        15'h2D7F: data = 12'h468;
        15'h2D80: data = 12'h453;
        15'h2D81: data = 12'h43F;
        15'h2D82: data = 12'h42C;
        15'h2D83: data = 12'h417;
        15'h2D84: data = 12'h402;
        15'h2D85: data = 12'h3E8;
        15'h2D86: data = 12'h3D2;
        15'h2D87: data = 12'h3C0;
        15'h2D88: data = 12'h3AE;
        15'h2D89: data = 12'h393;
        15'h2D8A: data = 12'h386;
        15'h2D8B: data = 12'h36F;
        15'h2D8C: data = 12'h358;
        15'h2D8D: data = 12'h345;
        15'h2D8E: data = 12'h32F;
        15'h2D8F: data = 12'h31D;
        15'h2D90: data = 12'h301;
        15'h2D91: data = 12'h2F1;
        15'h2D92: data = 12'h2D6;
        15'h2D93: data = 12'h2C4;
        15'h2D94: data = 12'h2A8;
        15'h2D95: data = 12'h290;
        15'h2D96: data = 12'h280;
        15'h2D97: data = 12'h265;
        15'h2D98: data = 12'h24D;
        15'h2D99: data = 12'h237;
        15'h2D9A: data = 12'h21E;
        15'h2D9B: data = 12'h208;
        15'h2D9C: data = 12'h1F7;
        15'h2D9D: data = 12'h1D8;
        15'h2D9E: data = 12'h1C1;
        15'h2D9F: data = 12'h1AA;
        15'h2DA0: data = 12'h192;
        15'h2DA1: data = 12'h17B;
        15'h2DA2: data = 12'h169;
        15'h2DA3: data = 12'h14F;
        15'h2DA4: data = 12'h139;
        15'h2DA5: data = 12'h11E;
        15'h2DA6: data = 12'h10A;
        15'h2DA7: data = 12'h0F5;
        15'h2DA8: data = 12'h0DB;
        15'h2DA9: data = 12'h0C0;
        15'h2DAA: data = 12'h0A8;
        15'h2DAB: data = 12'h091;
        15'h2DAC: data = 12'h07C;
        15'h2DAD: data = 12'h065;
        15'h2DAE: data = 12'h04E;
        15'h2DAF: data = 12'h7DF;
        15'h2DB0: data = 12'h7CE;
        15'h2DB1: data = 12'h7BD;
        15'h2DB2: data = 12'h7A3;
        15'h2DB3: data = 12'h78E;
        15'h2DB4: data = 12'h774;
        15'h2DB5: data = 12'h75C;
        15'h2DB6: data = 12'h749;
        15'h2DB7: data = 12'h732;
        15'h2DB8: data = 12'h71C;
        15'h2DB9: data = 12'h704;
        15'h2DBA: data = 12'h6EC;
        15'h2DBB: data = 12'h6D7;
        15'h2DBC: data = 12'h6C4;
        15'h2DBD: data = 12'h6AC;
        15'h2DBE: data = 12'h697;
        15'h2DBF: data = 12'h682;
        15'h2DC0: data = 12'h669;
        15'h2DC1: data = 12'h655;
        15'h2DC2: data = 12'h63B;
        15'h2DC3: data = 12'h62A;
        15'h2DC4: data = 12'h611;
        15'h2DC5: data = 12'h5F7;
        15'h2DC6: data = 12'h5DE;
        15'h2DC7: data = 12'h5CA;
        15'h2DC8: data = 12'h5B5;
        15'h2DC9: data = 12'h59C;
        15'h2DCA: data = 12'h584;
        15'h2DCB: data = 12'h56E;
        15'h2DCC: data = 12'h55C;
        15'h2DCD: data = 12'h546;
        15'h2DCE: data = 12'h533;
        15'h2DCF: data = 12'h51A;
        15'h2DD0: data = 12'h507;
        15'h2DD1: data = 12'h4F0;
        15'h2DD2: data = 12'h4DD;
        15'h2DD3: data = 12'h4CB;
        15'h2DD4: data = 12'h4B8;
        15'h2DD5: data = 12'h4A2;
        15'h2DD6: data = 12'h491;
        15'h2DD7: data = 12'h47C;
        15'h2DD8: data = 12'h46C;
        15'h2DD9: data = 12'h459;
        15'h2DDA: data = 12'h44D;
        15'h2DDB: data = 12'h43B;
        15'h2DDC: data = 12'h42C;
        15'h2DDD: data = 12'h419;
        15'h2DDE: data = 12'h408;
        15'h2DDF: data = 12'h3F6;
        15'h2DE0: data = 12'h3E7;
        15'h2DE1: data = 12'h3D2;
        15'h2DE2: data = 12'h3BE;
        15'h2DE3: data = 12'h3AF;
        15'h2DE4: data = 12'h399;
        15'h2DE5: data = 12'h391;
        15'h2DE6: data = 12'h376;
        15'h2DE7: data = 12'h362;
        15'h2DE8: data = 12'h350;
        15'h2DE9: data = 12'h33F;
        15'h2DEA: data = 12'h32E;
        15'h2DEB: data = 12'h31C;
        15'h2DEC: data = 12'h30C;
        15'h2DED: data = 12'h2FE;
        15'h2DEE: data = 12'h2F0;
        15'h2DEF: data = 12'h2E1;
        15'h2DF0: data = 12'h2D7;
        15'h2DF1: data = 12'h2D3;
        15'h2DF2: data = 12'h2C6;
        15'h2DF3: data = 12'h2B8;
        15'h2DF4: data = 12'h2AE;
        15'h2DF5: data = 12'h29F;
        15'h2DF6: data = 12'h296;
        15'h2DF7: data = 12'h283;
        15'h2DF8: data = 12'h27B;
        15'h2DF9: data = 12'h266;
        15'h2DFA: data = 12'h258;
        15'h2DFB: data = 12'h24A;
        15'h2DFC: data = 12'h23B;
        15'h2DFD: data = 12'h22D;
        15'h2DFE: data = 12'h221;
        15'h2DFF: data = 12'h216;
        15'h2E00: data = 12'h211;
        15'h2E01: data = 12'h20B;
        15'h2E02: data = 12'h20A;
        15'h2E03: data = 12'h1FC;
        15'h2E04: data = 12'h1F6;
        15'h2E05: data = 12'h1F0;
        15'h2E06: data = 12'h1E8;
        15'h2E07: data = 12'h1E0;
        15'h2E08: data = 12'h1D5;
        15'h2E09: data = 12'h1C8;
        15'h2E0A: data = 12'h1BC;
        15'h2E0B: data = 12'h1B9;
        15'h2E0C: data = 12'h1AC;
        15'h2E0D: data = 12'h1A3;
        15'h2E0E: data = 12'h19C;
        15'h2E0F: data = 12'h194;
        15'h2E10: data = 12'h190;
        15'h2E11: data = 12'h18E;
        15'h2E12: data = 12'h18A;
        15'h2E13: data = 12'h18A;
        15'h2E14: data = 12'h18D;
        15'h2E15: data = 12'h184;
        15'h2E16: data = 12'h186;
        15'h2E17: data = 12'h17E;
        15'h2E18: data = 12'h17F;
        15'h2E19: data = 12'h173;
        15'h2E1A: data = 12'h16F;
        15'h2E1B: data = 12'h16C;
        15'h2E1C: data = 12'h15C;
        15'h2E1D: data = 12'h160;
        15'h2E1E: data = 12'h15E;
        15'h2E1F: data = 12'h15E;
        15'h2E20: data = 12'h158;
        15'h2E21: data = 12'h159;
        15'h2E22: data = 12'h161;
        15'h2E23: data = 12'h164;
        15'h2E24: data = 12'h168;
        15'h2E25: data = 12'h169;
        15'h2E26: data = 12'h167;
        15'h2E27: data = 12'h170;
        15'h2E28: data = 12'h16E;
        15'h2E29: data = 12'h16E;
        15'h2E2A: data = 12'h168;
        15'h2E2B: data = 12'h164;
        15'h2E2C: data = 12'h166;
        15'h2E2D: data = 12'h163;
        15'h2E2E: data = 12'h169;
        15'h2E2F: data = 12'h169;
        15'h2E30: data = 12'h16E;
        15'h2E31: data = 12'h177;
        15'h2E32: data = 12'h182;
        15'h2E33: data = 12'h188;
        15'h2E34: data = 12'h191;
        15'h2E35: data = 12'h197;
        15'h2E36: data = 12'h19D;
        15'h2E37: data = 12'h1A5;
        15'h2E38: data = 12'h1AC;
        15'h2E39: data = 12'h1B3;
        15'h2E3A: data = 12'h1B2;
        15'h2E3B: data = 12'h1B3;
        15'h2E3C: data = 12'h1B6;
        15'h2E3D: data = 12'h1BA;
        15'h2E3E: data = 12'h1C2;
        15'h2E3F: data = 12'h1C6;
        15'h2E40: data = 12'h1CF;
        15'h2E41: data = 12'h1D8;
        15'h2E42: data = 12'h1E5;
        15'h2E43: data = 12'h1F3;
        15'h2E44: data = 12'h203;
        15'h2E45: data = 12'h20D;
        15'h2E46: data = 12'h21E;
        15'h2E47: data = 12'h220;
        15'h2E48: data = 12'h230;
        15'h2E49: data = 12'h237;
        15'h2E4A: data = 12'h246;
        15'h2E4B: data = 12'h24C;
        15'h2E4C: data = 12'h257;
        15'h2E4D: data = 12'h261;
        15'h2E4E: data = 12'h26B;
        15'h2E4F: data = 12'h26F;
        15'h2E50: data = 12'h279;
        15'h2E51: data = 12'h284;
        15'h2E52: data = 12'h291;
        15'h2E53: data = 12'h2A3;
        15'h2E54: data = 12'h2B3;
        15'h2E55: data = 12'h2C5;
        15'h2E56: data = 12'h2D3;
        15'h2E57: data = 12'h2E2;
        15'h2E58: data = 12'h2F5;
        15'h2E59: data = 12'h308;
        15'h2E5A: data = 12'h318;
        15'h2E5B: data = 12'h32A;
        15'h2E5C: data = 12'h335;
        15'h2E5D: data = 12'h344;
        15'h2E5E: data = 12'h352;
        15'h2E5F: data = 12'h360;
        15'h2E60: data = 12'h370;
        15'h2E61: data = 12'h37C;
        15'h2E62: data = 12'h38E;
        15'h2E63: data = 12'h393;
        15'h2E64: data = 12'h3A9;
        15'h2E65: data = 12'h3B9;
        15'h2E66: data = 12'h3C5;
        15'h2E67: data = 12'h3E0;
        15'h2E68: data = 12'h3EE;
        15'h2E69: data = 12'h400;
        15'h2E6A: data = 12'h419;
        15'h2E6B: data = 12'h42E;
        15'h2E6C: data = 12'h442;
        15'h2E6D: data = 12'h455;
        15'h2E6E: data = 12'h46A;
        15'h2E6F: data = 12'h485;
        15'h2E70: data = 12'h493;
        15'h2E71: data = 12'h4A8;
        15'h2E72: data = 12'h4B9;
        15'h2E73: data = 12'h4D0;
        15'h2E74: data = 12'h4E3;
        15'h2E75: data = 12'h4F4;
        15'h2E76: data = 12'h50A;
        15'h2E77: data = 12'h516;
        15'h2E78: data = 12'h525;
        15'h2E79: data = 12'h53C;
        15'h2E7A: data = 12'h551;
        15'h2E7B: data = 12'h564;
        15'h2E7C: data = 12'h573;
        15'h2E7D: data = 12'h589;
        15'h2E7E: data = 12'h5A2;
        15'h2E7F: data = 12'h5B9;
        15'h2E80: data = 12'h5CC;
        15'h2E81: data = 12'h5E7;
        15'h2E82: data = 12'h602;
        15'h2E83: data = 12'h61B;
        15'h2E84: data = 12'h631;
        15'h2E85: data = 12'h648;
        15'h2E86: data = 12'h664;
        15'h2E87: data = 12'h677;
        15'h2E88: data = 12'h692;
        15'h2E89: data = 12'h6A4;
        15'h2E8A: data = 12'h6B9;
        15'h2E8B: data = 12'h6CD;
        15'h2E8C: data = 12'h6E0;
        15'h2E8D: data = 12'h6F3;
        15'h2E8E: data = 12'h708;
        15'h2E8F: data = 12'h71C;
        15'h2E90: data = 12'h734;
        15'h2E91: data = 12'h745;
        15'h2E92: data = 12'h75B;
        15'h2E93: data = 12'h775;
        15'h2E94: data = 12'h791;
        15'h2E95: data = 12'h79F;
        15'h2E96: data = 12'h7B8;
        15'h2E97: data = 12'h7D6;
        15'h2E98: data = 12'h7ED;
        15'h2E99: data = 12'h804;
        15'h2E9A: data = 12'h077;
        15'h2E9B: data = 12'h08D;
        15'h2E9C: data = 12'h0A3;
        15'h2E9D: data = 12'h0B5;
        15'h2E9E: data = 12'h0D1;
        15'h2E9F: data = 12'h0EA;
        15'h2EA0: data = 12'h102;
        15'h2EA1: data = 12'h112;
        15'h2EA2: data = 12'h12A;
        15'h2EA3: data = 12'h144;
        15'h2EA4: data = 12'h155;
        15'h2EA5: data = 12'h16B;
        15'h2EA6: data = 12'h17E;
        15'h2EA7: data = 12'h199;
        15'h2EA8: data = 12'h1AE;
        15'h2EA9: data = 12'h1BD;
        15'h2EAA: data = 12'h1D5;
        15'h2EAB: data = 12'h1ED;
        15'h2EAC: data = 12'h204;
        15'h2EAD: data = 12'h218;
        15'h2EAE: data = 12'h231;
        15'h2EAF: data = 12'h24A;
        15'h2EB0: data = 12'h263;
        15'h2EB1: data = 12'h275;
        15'h2EB2: data = 12'h28C;
        15'h2EB3: data = 12'h2A8;
        15'h2EB4: data = 12'h2C3;
        15'h2EB5: data = 12'h2D8;
        15'h2EB6: data = 12'h2F4;
        15'h2EB7: data = 12'h30D;
        15'h2EB8: data = 12'h327;
        15'h2EB9: data = 12'h338;
        15'h2EBA: data = 12'h34D;
        15'h2EBB: data = 12'h368;
        15'h2EBC: data = 12'h380;
        15'h2EBD: data = 12'h398;
        15'h2EBE: data = 12'h3AB;
        15'h2EBF: data = 12'h3C8;
        15'h2EC0: data = 12'h3DD;
        15'h2EC1: data = 12'h3F2;
        15'h2EC2: data = 12'h3FF;
        15'h2EC3: data = 12'h417;
        15'h2EC4: data = 12'h42E;
        15'h2EC5: data = 12'h446;
        15'h2EC6: data = 12'h455;
        15'h2EC7: data = 12'h469;
        15'h2EC8: data = 12'h47F;
        15'h2EC9: data = 12'h492;
        15'h2ECA: data = 12'h4A6;
        15'h2ECB: data = 12'h4B9;
        15'h2ECC: data = 12'h4C5;
        15'h2ECD: data = 12'h4D8;
        15'h2ECE: data = 12'h4EE;
        15'h2ECF: data = 12'h503;
        15'h2ED0: data = 12'h510;
        15'h2ED1: data = 12'h526;
        15'h2ED2: data = 12'h53B;
        15'h2ED3: data = 12'h54B;
        15'h2ED4: data = 12'h55B;
        15'h2ED5: data = 12'h569;
        15'h2ED6: data = 12'h582;
        15'h2ED7: data = 12'h593;
        15'h2ED8: data = 12'h5A7;
        15'h2ED9: data = 12'h5BB;
        15'h2EDA: data = 12'h5C2;
        15'h2EDB: data = 12'h5DB;
        15'h2EDC: data = 12'h5EE;
        15'h2EDD: data = 12'h5FC;
        15'h2EDE: data = 12'h60A;
        15'h2EDF: data = 12'h61B;
        15'h2EE0: data = 12'h62C;
        15'h2EE1: data = 12'h63D;
        15'h2EE2: data = 12'h654;
        15'h2EE3: data = 12'h665;
        15'h2EE4: data = 12'h676;
        15'h2EE5: data = 12'h683;
        15'h2EE6: data = 12'h694;
        15'h2EE7: data = 12'h6A2;
        15'h2EE8: data = 12'h6B2;
        15'h2EE9: data = 12'h6C1;
        15'h2EEA: data = 12'h6D3;
        15'h2EEB: data = 12'h6DD;
        15'h2EEC: data = 12'h6ED;
        15'h2EED: data = 12'h6FD;
        15'h2EEE: data = 12'h707;
        15'h2EEF: data = 12'h710;
        15'h2EF0: data = 12'h724;
        15'h2EF1: data = 12'h732;
        15'h2EF2: data = 12'h73C;
        15'h2EF3: data = 12'h744;
        15'h2EF4: data = 12'h74E;
        15'h2EF5: data = 12'h760;
        15'h2EF6: data = 12'h768;
        15'h2EF7: data = 12'h778;
        15'h2EF8: data = 12'h77B;
        15'h2EF9: data = 12'h78D;
        15'h2EFA: data = 12'h795;
        15'h2EFB: data = 12'h79C;
        15'h2EFC: data = 12'h7A4;
        15'h2EFD: data = 12'h7AF;
        15'h2EFE: data = 12'h7B9;
        15'h2EFF: data = 12'h7BD;
        15'h2F00: data = 12'h7C7;
        15'h2F01: data = 12'h7CE;
        15'h2F02: data = 12'h7D6;
        15'h2F03: data = 12'h7DB;
        15'h2F04: data = 12'h7E9;
        15'h2F05: data = 12'h7EE;
        15'h2F06: data = 12'h7F1;
        15'h2F07: data = 12'h7F8;
        15'h2F08: data = 12'h801;
        15'h2F09: data = 12'h803;
        15'h2F0A: data = 12'h805;
        15'h2F0B: data = 12'h80D;
        15'h2F0C: data = 12'h07B;
        15'h2F0D: data = 12'h08A;
        15'h2F0E: data = 12'h095;
        15'h2F0F: data = 12'h09A;
        15'h2F10: data = 12'h098;
        15'h2F11: data = 12'h09E;
        15'h2F12: data = 12'h0A0;
        15'h2F13: data = 12'h0AB;
        15'h2F14: data = 12'h0AB;
        15'h2F15: data = 12'h0AE;
        15'h2F16: data = 12'h0B4;
        15'h2F17: data = 12'h0B9;
        15'h2F18: data = 12'h0BA;
        15'h2F19: data = 12'h0B8;
        15'h2F1A: data = 12'h0C5;
        15'h2F1B: data = 12'h0C9;
        15'h2F1C: data = 12'h0C9;
        15'h2F1D: data = 12'h0CF;
        15'h2F1E: data = 12'h0D3;
        15'h2F1F: data = 12'h0D2;
        15'h2F20: data = 12'h0D4;
        15'h2F21: data = 12'h0D0;
        15'h2F22: data = 12'h0D0;
        15'h2F23: data = 12'h0CC;
        15'h2F24: data = 12'h0CD;
        15'h2F25: data = 12'h0C5;
        15'h2F26: data = 12'h0BD;
        15'h2F27: data = 12'h0B9;
        15'h2F28: data = 12'h0B0;
        15'h2F29: data = 12'h0AF;
        15'h2F2A: data = 12'h0A6;
        15'h2F2B: data = 12'h0A8;
        15'h2F2C: data = 12'h0AC;
        15'h2F2D: data = 12'h0B0;
        15'h2F2E: data = 12'h0AC;
        15'h2F2F: data = 12'h0A7;
        15'h2F30: data = 12'h0A6;
        15'h2F31: data = 12'h09B;
        15'h2F32: data = 12'h090;
        15'h2F33: data = 12'h083;
        15'h2F34: data = 12'h077;
        15'h2F35: data = 12'h076;
        15'h2F36: data = 12'h06F;
        15'h2F37: data = 12'h06B;
        15'h2F38: data = 12'h06B;
        15'h2F39: data = 12'h068;
        15'h2F3A: data = 12'h05F;
        15'h2F3B: data = 12'h057;
        15'h2F3C: data = 12'h045;
        15'h2F3D: data = 12'h7C0;
        15'h2F3E: data = 12'h7B4;
        15'h2F3F: data = 12'h7A7;
        15'h2F40: data = 12'h7A1;
        15'h2F41: data = 12'h793;
        15'h2F42: data = 12'h794;
        15'h2F43: data = 12'h78A;
        15'h2F44: data = 12'h77D;
        15'h2F45: data = 12'h76B;
        15'h2F46: data = 12'h759;
        15'h2F47: data = 12'h744;
        15'h2F48: data = 12'h736;
        15'h2F49: data = 12'h72D;
        15'h2F4A: data = 12'h727;
        15'h2F4B: data = 12'h71B;
        15'h2F4C: data = 12'h711;
        15'h2F4D: data = 12'h70A;
        15'h2F4E: data = 12'h6FB;
        15'h2F4F: data = 12'h6EB;
        15'h2F50: data = 12'h6DD;
        15'h2F51: data = 12'h6CC;
        15'h2F52: data = 12'h6B4;
        15'h2F53: data = 12'h6A3;
        15'h2F54: data = 12'h693;
        15'h2F55: data = 12'h687;
        15'h2F56: data = 12'h67E;
        15'h2F57: data = 12'h671;
        15'h2F58: data = 12'h667;
        15'h2F59: data = 12'h656;
        15'h2F5A: data = 12'h646;
        15'h2F5B: data = 12'h635;
        15'h2F5C: data = 12'h62A;
        15'h2F5D: data = 12'h611;
        15'h2F5E: data = 12'h5FC;
        15'h2F5F: data = 12'h5EA;
        15'h2F60: data = 12'h5D0;
        15'h2F61: data = 12'h5BF;
        15'h2F62: data = 12'h5AE;
        15'h2F63: data = 12'h5A2;
        15'h2F64: data = 12'h58E;
        15'h2F65: data = 12'h57D;
        15'h2F66: data = 12'h56F;
        15'h2F67: data = 12'h563;
        15'h2F68: data = 12'h558;
        15'h2F69: data = 12'h546;
        15'h2F6A: data = 12'h52D;
        15'h2F6B: data = 12'h519;
        15'h2F6C: data = 12'h506;
        15'h2F6D: data = 12'h4F1;
        15'h2F6E: data = 12'h4DB;
        15'h2F6F: data = 12'h4C1;
        15'h2F70: data = 12'h4AF;
        15'h2F71: data = 12'h498;
        15'h2F72: data = 12'h480;
        15'h2F73: data = 12'h469;
        15'h2F74: data = 12'h452;
        15'h2F75: data = 12'h441;
        15'h2F76: data = 12'h42B;
        15'h2F77: data = 12'h412;
        15'h2F78: data = 12'h3FF;
        15'h2F79: data = 12'h3E7;
        15'h2F7A: data = 12'h3D0;
        15'h2F7B: data = 12'h3BF;
        15'h2F7C: data = 12'h3AC;
        15'h2F7D: data = 12'h392;
        15'h2F7E: data = 12'h37F;
        15'h2F7F: data = 12'h369;
        15'h2F80: data = 12'h352;
        15'h2F81: data = 12'h340;
        15'h2F82: data = 12'h32D;
        15'h2F83: data = 12'h318;
        15'h2F84: data = 12'h2FE;
        15'h2F85: data = 12'h2EA;
        15'h2F86: data = 12'h2D7;
        15'h2F87: data = 12'h2BF;
        15'h2F88: data = 12'h2A7;
        15'h2F89: data = 12'h290;
        15'h2F8A: data = 12'h27C;
        15'h2F8B: data = 12'h268;
        15'h2F8C: data = 12'h24C;
        15'h2F8D: data = 12'h236;
        15'h2F8E: data = 12'h21A;
        15'h2F8F: data = 12'h209;
        15'h2F90: data = 12'h1F3;
        15'h2F91: data = 12'h1DA;
        15'h2F92: data = 12'h1BF;
        15'h2F93: data = 12'h1A9;
        15'h2F94: data = 12'h192;
        15'h2F95: data = 12'h17F;
        15'h2F96: data = 12'h169;
        15'h2F97: data = 12'h153;
        15'h2F98: data = 12'h13A;
        15'h2F99: data = 12'h11F;
        15'h2F9A: data = 12'h109;
        15'h2F9B: data = 12'h0F2;
        15'h2F9C: data = 12'h0DC;
        15'h2F9D: data = 12'h0C2;
        15'h2F9E: data = 12'h0A9;
        15'h2F9F: data = 12'h092;
        15'h2FA0: data = 12'h080;
        15'h2FA1: data = 12'h067;
        15'h2FA2: data = 12'h050;
        15'h2FA3: data = 12'h7E1;
        15'h2FA4: data = 12'h7CD;
        15'h2FA5: data = 12'h7BD;
        15'h2FA6: data = 12'h7A3;
        15'h2FA7: data = 12'h78C;
        15'h2FA8: data = 12'h779;
        15'h2FA9: data = 12'h75C;
        15'h2FAA: data = 12'h74B;
        15'h2FAB: data = 12'h734;
        15'h2FAC: data = 12'h722;
        15'h2FAD: data = 12'h708;
        15'h2FAE: data = 12'h6E9;
        15'h2FAF: data = 12'h6D7;
        15'h2FB0: data = 12'h6C3;
        15'h2FB1: data = 12'h6AD;
        15'h2FB2: data = 12'h697;
        15'h2FB3: data = 12'h681;
        15'h2FB4: data = 12'h668;
        15'h2FB5: data = 12'h656;
        15'h2FB6: data = 12'h63D;
        15'h2FB7: data = 12'h62D;
        15'h2FB8: data = 12'h615;
        15'h2FB9: data = 12'h5FB;
        15'h2FBA: data = 12'h5E6;
        15'h2FBB: data = 12'h5D0;
        15'h2FBC: data = 12'h5BB;
        15'h2FBD: data = 12'h59E;
        15'h2FBE: data = 12'h587;
        15'h2FBF: data = 12'h575;
        15'h2FC0: data = 12'h560;
        15'h2FC1: data = 12'h549;
        15'h2FC2: data = 12'h538;
        15'h2FC3: data = 12'h51E;
        15'h2FC4: data = 12'h50A;
        15'h2FC5: data = 12'h4F4;
        15'h2FC6: data = 12'h4DF;
        15'h2FC7: data = 12'h4CD;
        15'h2FC8: data = 12'h4B8;
        15'h2FC9: data = 12'h4A2;
        15'h2FCA: data = 12'h48F;
        15'h2FCB: data = 12'h47E;
        15'h2FCC: data = 12'h468;
        15'h2FCD: data = 12'h45A;
        15'h2FCE: data = 12'h44D;
        15'h2FCF: data = 12'h43A;
        15'h2FD0: data = 12'h429;
        15'h2FD1: data = 12'h416;
        15'h2FD2: data = 12'h402;
        15'h2FD3: data = 12'h3F5;
        15'h2FD4: data = 12'h3E7;
        15'h2FD5: data = 12'h3D0;
        15'h2FD6: data = 12'h3C3;
        15'h2FD7: data = 12'h3AF;
        15'h2FD8: data = 12'h39F;
        15'h2FD9: data = 12'h392;
        15'h2FDA: data = 12'h378;
        15'h2FDB: data = 12'h364;
        15'h2FDC: data = 12'h354;
        15'h2FDD: data = 12'h341;
        15'h2FDE: data = 12'h330;
        15'h2FDF: data = 12'h31F;
        15'h2FE0: data = 12'h310;
        15'h2FE1: data = 12'h300;
        15'h2FE2: data = 12'h2F1;
        15'h2FE3: data = 12'h2E3;
        15'h2FE4: data = 12'h2D4;
        15'h2FE5: data = 12'h2D2;
        15'h2FE6: data = 12'h2C7;
        15'h2FE7: data = 12'h2B9;
        15'h2FE8: data = 12'h2AB;
        15'h2FE9: data = 12'h2A2;
        15'h2FEA: data = 12'h293;
        15'h2FEB: data = 12'h283;
        15'h2FEC: data = 12'h27C;
        15'h2FED: data = 12'h269;
        15'h2FEE: data = 12'h260;
        15'h2FEF: data = 12'h24D;
        15'h2FF0: data = 12'h240;
        15'h2FF1: data = 12'h230;
        15'h2FF2: data = 12'h224;
        15'h2FF3: data = 12'h217;
        15'h2FF4: data = 12'h20E;
        15'h2FF5: data = 12'h209;
        15'h2FF6: data = 12'h204;
        15'h2FF7: data = 12'h1F7;
        15'h2FF8: data = 12'h1F6;
        15'h2FF9: data = 12'h1F1;
        15'h2FFA: data = 12'h1EE;
        15'h2FFB: data = 12'h1E3;
        15'h2FFC: data = 12'h1D7;
        15'h2FFD: data = 12'h1CA;
        15'h2FFE: data = 12'h1C3;
        15'h2FFF: data = 12'h1BD;
        15'h3000: data = 12'h1B0;
        15'h3001: data = 12'h1A6;
        15'h3002: data = 12'h19B;
        15'h3003: data = 12'h194;
        15'h3004: data = 12'h191;
        15'h3005: data = 12'h18C;
        15'h3006: data = 12'h187;
        15'h3007: data = 12'h186;
        15'h3008: data = 12'h18B;
        15'h3009: data = 12'h180;
        15'h300A: data = 12'h185;
        15'h300B: data = 12'h17D;
        15'h300C: data = 12'h17E;
        15'h300D: data = 12'h174;
        15'h300E: data = 12'h173;
        15'h300F: data = 12'h170;
        15'h3010: data = 12'h161;
        15'h3011: data = 12'h160;
        15'h3012: data = 12'h15B;
        15'h3013: data = 12'h15A;
        15'h3014: data = 12'h156;
        15'h3015: data = 12'h15B;
        15'h3016: data = 12'h15D;
        15'h3017: data = 12'h161;
        15'h3018: data = 12'h166;
        15'h3019: data = 12'h165;
        15'h301A: data = 12'h167;
        15'h301B: data = 12'h16E;
        15'h301C: data = 12'h16C;
        15'h301D: data = 12'h16D;
        15'h301E: data = 12'h16A;
        15'h301F: data = 12'h165;
        15'h3020: data = 12'h16A;
        15'h3021: data = 12'h169;
        15'h3022: data = 12'h168;
        15'h3023: data = 12'h16D;
        15'h3024: data = 12'h16A;
        15'h3025: data = 12'h175;
        15'h3026: data = 12'h182;
        15'h3027: data = 12'h185;
        15'h3028: data = 12'h192;
        15'h3029: data = 12'h193;
        15'h302A: data = 12'h19A;
        15'h302B: data = 12'h1A4;
        15'h302C: data = 12'h1AB;
        15'h302D: data = 12'h1B1;
        15'h302E: data = 12'h1B3;
        15'h302F: data = 12'h1B6;
        15'h3030: data = 12'h1B8;
        15'h3031: data = 12'h1BC;
        15'h3032: data = 12'h1C0;
        15'h3033: data = 12'h1C9;
        15'h3034: data = 12'h1D0;
        15'h3035: data = 12'h1D6;
        15'h3036: data = 12'h1E2;
        15'h3037: data = 12'h1F0;
        15'h3038: data = 12'h1FE;
        15'h3039: data = 12'h208;
        15'h303A: data = 12'h218;
        15'h303B: data = 12'h21D;
        15'h303C: data = 12'h22D;
        15'h303D: data = 12'h238;
        15'h303E: data = 12'h246;
        15'h303F: data = 12'h24F;
        15'h3040: data = 12'h25B;
        15'h3041: data = 12'h265;
        15'h3042: data = 12'h26B;
        15'h3043: data = 12'h273;
        15'h3044: data = 12'h27E;
        15'h3045: data = 12'h289;
        15'h3046: data = 12'h292;
        15'h3047: data = 12'h2A1;
        15'h3048: data = 12'h2B2;
        15'h3049: data = 12'h2C0;
        15'h304A: data = 12'h2D0;
        15'h304B: data = 12'h2DE;
        15'h304C: data = 12'h2F2;
        15'h304D: data = 12'h306;
        15'h304E: data = 12'h313;
        15'h304F: data = 12'h326;
        15'h3050: data = 12'h339;
        15'h3051: data = 12'h346;
        15'h3052: data = 12'h355;
        15'h3053: data = 12'h366;
        15'h3054: data = 12'h36F;
        15'h3055: data = 12'h381;
        15'h3056: data = 12'h392;
        15'h3057: data = 12'h398;
        15'h3058: data = 12'h3AA;
        15'h3059: data = 12'h3B7;
        15'h305A: data = 12'h3C6;
        15'h305B: data = 12'h3DC;
        15'h305C: data = 12'h3EA;
        15'h305D: data = 12'h3FC;
        15'h305E: data = 12'h416;
        15'h305F: data = 12'h42A;
        15'h3060: data = 12'h440;
        15'h3061: data = 12'h451;
        15'h3062: data = 12'h466;
        15'h3063: data = 12'h484;
        15'h3064: data = 12'h494;
        15'h3065: data = 12'h4A8;
        15'h3066: data = 12'h4B7;
        15'h3067: data = 12'h4CE;
        15'h3068: data = 12'h4E2;
        15'h3069: data = 12'h4F7;
        15'h306A: data = 12'h50B;
        15'h306B: data = 12'h51C;
        15'h306C: data = 12'h52B;
        15'h306D: data = 12'h541;
        15'h306E: data = 12'h554;
        15'h306F: data = 12'h566;
        15'h3070: data = 12'h572;
        15'h3071: data = 12'h589;
        15'h3072: data = 12'h59F;
        15'h3073: data = 12'h5B6;
        15'h3074: data = 12'h5CA;
        15'h3075: data = 12'h5E5;
        15'h3076: data = 12'h5FC;
        15'h3077: data = 12'h616;
        15'h3078: data = 12'h62D;
        15'h3079: data = 12'h645;
        15'h307A: data = 12'h660;
        15'h307B: data = 12'h678;
        15'h307C: data = 12'h690;
        15'h307D: data = 12'h6A1;
        15'h307E: data = 12'h6B7;
        15'h307F: data = 12'h6CE;
        15'h3080: data = 12'h6E3;
        15'h3081: data = 12'h6F5;
        15'h3082: data = 12'h70E;
        15'h3083: data = 12'h722;
        15'h3084: data = 12'h736;
        15'h3085: data = 12'h745;
        15'h3086: data = 12'h75A;
        15'h3087: data = 12'h775;
        15'h3088: data = 12'h78D;
        15'h3089: data = 12'h79D;
        15'h308A: data = 12'h7B7;
        15'h308B: data = 12'h7D0;
        15'h308C: data = 12'h7E8;
        15'h308D: data = 12'h801;
        15'h308E: data = 12'h070;
        15'h308F: data = 12'h088;
        15'h3090: data = 12'h09E;
        15'h3091: data = 12'h0B3;
        15'h3092: data = 12'h0CF;
        15'h3093: data = 12'h0E6;
        15'h3094: data = 12'h0FE;
        15'h3095: data = 12'h113;
        15'h3096: data = 12'h12C;
        15'h3097: data = 12'h146;
        15'h3098: data = 12'h15B;
        15'h3099: data = 12'h16F;
        15'h309A: data = 12'h183;
        15'h309B: data = 12'h19C;
        15'h309C: data = 12'h1B5;
        15'h309D: data = 12'h1C2;
        15'h309E: data = 12'h1D9;
        15'h309F: data = 12'h1EE;
        15'h30A0: data = 12'h206;
        15'h30A1: data = 12'h21A;
        15'h30A2: data = 12'h232;
        15'h30A3: data = 12'h24C;
        15'h30A4: data = 12'h264;
        15'h30A5: data = 12'h277;
        15'h30A6: data = 12'h28B;
        15'h30A7: data = 12'h2A6;
        15'h30A8: data = 12'h2BE;
        15'h30A9: data = 12'h2D1;
        15'h30AA: data = 12'h2EE;
        15'h30AB: data = 12'h306;
        15'h30AC: data = 12'h322;
        15'h30AD: data = 12'h334;
        15'h30AE: data = 12'h34D;
        15'h30AF: data = 12'h366;
        15'h30B0: data = 12'h37E;
        15'h30B1: data = 12'h397;
        15'h30B2: data = 12'h3AC;
        15'h30B3: data = 12'h3C5;
        15'h30B4: data = 12'h3DE;
        15'h30B5: data = 12'h3F2;
        15'h30B6: data = 12'h3FE;
        15'h30B7: data = 12'h417;
        15'h30B8: data = 12'h42C;
        15'h30B9: data = 12'h445;
        15'h30BA: data = 12'h452;
        15'h30BB: data = 12'h467;
        15'h30BC: data = 12'h47E;
        15'h30BD: data = 12'h494;
        15'h30BE: data = 12'h4AB;
        15'h30BF: data = 12'h4B9;
        15'h30C0: data = 12'h4C9;
        15'h30C1: data = 12'h4DA;
        15'h30C2: data = 12'h4F1;
        15'h30C3: data = 12'h506;
        15'h30C4: data = 12'h513;
        15'h30C5: data = 12'h526;
        15'h30C6: data = 12'h53B;
        15'h30C7: data = 12'h54C;
        15'h30C8: data = 12'h55F;
        15'h30C9: data = 12'h56C;
        15'h30CA: data = 12'h582;
        15'h30CB: data = 12'h592;
        15'h30CC: data = 12'h5A8;
        15'h30CD: data = 12'h5B9;
        15'h30CE: data = 12'h5C8;
        15'h30CF: data = 12'h5D4;
        15'h30D0: data = 12'h5ED;
        15'h30D1: data = 12'h5FC;
        15'h30D2: data = 12'h60C;
        15'h30D3: data = 12'h61B;
        15'h30D4: data = 12'h627;
        15'h30D5: data = 12'h638;
        15'h30D6: data = 12'h650;
        15'h30D7: data = 12'h661;
        15'h30D8: data = 12'h672;
        15'h30D9: data = 12'h684;
        15'h30DA: data = 12'h696;
        15'h30DB: data = 12'h6A3;
        15'h30DC: data = 12'h6B3;
        15'h30DD: data = 12'h6C4;
        15'h30DE: data = 12'h6D2;
        15'h30DF: data = 12'h6DE;
        15'h30E0: data = 12'h6F0;
        15'h30E1: data = 12'h6FB;
        15'h30E2: data = 12'h709;
        15'h30E3: data = 12'h717;
        15'h30E4: data = 12'h726;
        15'h30E5: data = 12'h731;
        15'h30E6: data = 12'h73B;
        15'h30E7: data = 12'h74A;
        15'h30E8: data = 12'h74F;
        15'h30E9: data = 12'h761;
        15'h30EA: data = 12'h768;
        15'h30EB: data = 12'h775;
        15'h30EC: data = 12'h77E;
        15'h30ED: data = 12'h78E;
        15'h30EE: data = 12'h794;
        15'h30EF: data = 12'h79B;
        15'h30F0: data = 12'h7A2;
        15'h30F1: data = 12'h7AD;
        15'h30F2: data = 12'h7B6;
        15'h30F3: data = 12'h7BE;
        15'h30F4: data = 12'h7C8;
        15'h30F5: data = 12'h7CF;
        15'h30F6: data = 12'h7D6;
        15'h30F7: data = 12'h7DD;
        15'h30F8: data = 12'h7EA;
        15'h30F9: data = 12'h7EE;
        15'h30FA: data = 12'h7EF;
        15'h30FB: data = 12'h7F7;
        15'h30FC: data = 12'h7FE;
        15'h30FD: data = 12'h802;
        15'h30FE: data = 12'h801;
        15'h30FF: data = 12'h80A;
        15'h3100: data = 12'h78A;
        15'h3101: data = 12'h089;
        15'h3102: data = 12'h091;
        15'h3103: data = 12'h095;
        15'h3104: data = 12'h094;
        15'h3105: data = 12'h0A1;
        15'h3106: data = 12'h09F;
        15'h3107: data = 12'h0AA;
        15'h3108: data = 12'h0A7;
        15'h3109: data = 12'h0AC;
        15'h310A: data = 12'h0B4;
        15'h310B: data = 12'h0B8;
        15'h310C: data = 12'h0B9;
        15'h310D: data = 12'h0BA;
        15'h310E: data = 12'h0C8;
        15'h310F: data = 12'h0C9;
        15'h3110: data = 12'h0CF;
        15'h3111: data = 12'h0D3;
        15'h3112: data = 12'h0D1;
        15'h3113: data = 12'h0D2;
        15'h3114: data = 12'h0D5;
        15'h3115: data = 12'h0CE;
        15'h3116: data = 12'h0CC;
        15'h3117: data = 12'h0CC;
        15'h3118: data = 12'h0CA;
        15'h3119: data = 12'h0C4;
        15'h311A: data = 12'h0BC;
        15'h311B: data = 12'h0B5;
        15'h311C: data = 12'h0AC;
        15'h311D: data = 12'h0AC;
        15'h311E: data = 12'h0A7;
        15'h311F: data = 12'h0A8;
        15'h3120: data = 12'h0A9;
        15'h3121: data = 12'h0AF;
        15'h3122: data = 12'h0AD;
        15'h3123: data = 12'h0A5;
        15'h3124: data = 12'h0A4;
        15'h3125: data = 12'h09A;
        15'h3126: data = 12'h08D;
        15'h3127: data = 12'h080;
        15'h3128: data = 12'h074;
        15'h3129: data = 12'h073;
        15'h312A: data = 12'h06F;
        15'h312B: data = 12'h069;
        15'h312C: data = 12'h069;
        15'h312D: data = 12'h066;
        15'h312E: data = 12'h05F;
        15'h312F: data = 12'h053;
        15'h3130: data = 12'h043;
        15'h3131: data = 12'h7BF;
        15'h3132: data = 12'h7B4;
        15'h3133: data = 12'h7A5;
        15'h3134: data = 12'h7A1;
        15'h3135: data = 12'h798;
        15'h3136: data = 12'h792;
        15'h3137: data = 12'h78A;
        15'h3138: data = 12'h77C;
        15'h3139: data = 12'h768;
        15'h313A: data = 12'h758;
        15'h313B: data = 12'h745;
        15'h313C: data = 12'h738;
        15'h313D: data = 12'h72D;
        15'h313E: data = 12'h724;
        15'h313F: data = 12'h717;
        15'h3140: data = 12'h712;
        15'h3141: data = 12'h709;
        15'h3142: data = 12'h6FA;
        15'h3143: data = 12'h6EA;
        15'h3144: data = 12'h6DB;
        15'h3145: data = 12'h6C9;
        15'h3146: data = 12'h6B1;
        15'h3147: data = 12'h6A4;
        15'h3148: data = 12'h692;
        15'h3149: data = 12'h684;
        15'h314A: data = 12'h67A;
        15'h314B: data = 12'h66E;
        15'h314C: data = 12'h665;
        15'h314D: data = 12'h655;
        15'h314E: data = 12'h644;
        15'h314F: data = 12'h631;
        15'h3150: data = 12'h628;
        15'h3151: data = 12'h612;
        15'h3152: data = 12'h5FD;
        15'h3153: data = 12'h5E7;
        15'h3154: data = 12'h5CF;
        15'h3155: data = 12'h5BF;
        15'h3156: data = 12'h5B3;
        15'h3157: data = 12'h59F;
        15'h3158: data = 12'h58E;
        15'h3159: data = 12'h57C;
        15'h315A: data = 12'h56F;
        15'h315B: data = 12'h561;
        15'h315C: data = 12'h552;
        15'h315D: data = 12'h540;
        15'h315E: data = 12'h52B;
        15'h315F: data = 12'h518;
        15'h3160: data = 12'h503;
        15'h3161: data = 12'h4F4;
        15'h3162: data = 12'h4DC;
        15'h3163: data = 12'h4C7;
        15'h3164: data = 12'h4B3;
        15'h3165: data = 12'h499;
        15'h3166: data = 12'h482;
        15'h3167: data = 12'h46A;
        15'h3168: data = 12'h452;
        15'h3169: data = 12'h43D;
        15'h316A: data = 12'h42B;
        15'h316B: data = 12'h412;
        15'h316C: data = 12'h3FB;
        15'h316D: data = 12'h3E5;
        15'h316E: data = 12'h3D0;
        15'h316F: data = 12'h3BB;
        15'h3170: data = 12'h3A9;
        15'h3171: data = 12'h38F;
        15'h3172: data = 12'h37F;
        15'h3173: data = 12'h366;
        15'h3174: data = 12'h34F;
        15'h3175: data = 12'h33A;
        15'h3176: data = 12'h327;
        15'h3177: data = 12'h314;
        15'h3178: data = 12'h2FA;
        15'h3179: data = 12'h2E6;
        15'h317A: data = 12'h2D1;
        15'h317B: data = 12'h2BF;
        15'h317C: data = 12'h2A6;
        15'h317D: data = 12'h28D;
        15'h317E: data = 12'h27D;
        15'h317F: data = 12'h262;
        15'h3180: data = 12'h248;
        15'h3181: data = 12'h235;
        15'h3182: data = 12'h21C;
        15'h3183: data = 12'h201;
        15'h3184: data = 12'h1F4;
        15'h3185: data = 12'h1D6;
        15'h3186: data = 12'h1C1;
        15'h3187: data = 12'h1A9;
        15'h3188: data = 12'h192;
        15'h3189: data = 12'h17C;
        15'h318A: data = 12'h165;
        15'h318B: data = 12'h14F;
        15'h318C: data = 12'h136;
        15'h318D: data = 12'h121;
        15'h318E: data = 12'h109;
        15'h318F: data = 12'h0F3;
        15'h3190: data = 12'h0D9;
        15'h3191: data = 12'h0BE;
        15'h3192: data = 12'h0A8;
        15'h3193: data = 12'h08F;
        15'h3194: data = 12'h07F;
        15'h3195: data = 12'h063;
        15'h3196: data = 12'h04B;
        15'h3197: data = 12'h509;
        15'h3198: data = 12'h7CD;
        15'h3199: data = 12'h7BA;
        15'h319A: data = 12'h7A6;
        15'h319B: data = 12'h78F;
        15'h319C: data = 12'h776;
        15'h319D: data = 12'h75D;
        15'h319E: data = 12'h74B;
        15'h319F: data = 12'h734;
        15'h31A0: data = 12'h71C;
        15'h31A1: data = 12'h706;
        15'h31A2: data = 12'h6ED;
        15'h31A3: data = 12'h6D8;
        15'h31A4: data = 12'h6C3;
        15'h31A5: data = 12'h6AC;
        15'h31A6: data = 12'h695;
        15'h31A7: data = 12'h683;
        15'h31A8: data = 12'h668;
        15'h31A9: data = 12'h654;
        15'h31AA: data = 12'h63A;
        15'h31AB: data = 12'h62C;
        15'h31AC: data = 12'h614;
        15'h31AD: data = 12'h5FB;
        15'h31AE: data = 12'h5E4;
        15'h31AF: data = 12'h5CD;
        15'h31B0: data = 12'h5BA;
        15'h31B1: data = 12'h5A0;
        15'h31B2: data = 12'h58A;
        15'h31B3: data = 12'h574;
        15'h31B4: data = 12'h561;
        15'h31B5: data = 12'h54A;
        15'h31B6: data = 12'h535;
        15'h31B7: data = 12'h51E;
        15'h31B8: data = 12'h507;
        15'h31B9: data = 12'h4F5;
        15'h31BA: data = 12'h4DE;
        15'h31BB: data = 12'h4C7;
        15'h31BC: data = 12'h4B2;
        15'h31BD: data = 12'h4A2;
        15'h31BE: data = 12'h48F;
        15'h31BF: data = 12'h47A;
        15'h31C0: data = 12'h467;
        15'h31C1: data = 12'h457;
        15'h31C2: data = 12'h447;
        15'h31C3: data = 12'h437;
        15'h31C4: data = 12'h424;
        15'h31C5: data = 12'h413;
        15'h31C6: data = 12'h404;
        15'h31C7: data = 12'h3F8;
        15'h31C8: data = 12'h3E8;
        15'h31C9: data = 12'h3D0;
        15'h31CA: data = 12'h3C2;
        15'h31CB: data = 12'h3B0;
        15'h31CC: data = 12'h39E;
        15'h31CD: data = 12'h392;
        15'h31CE: data = 12'h37A;
        15'h31CF: data = 12'h36A;
        15'h31D0: data = 12'h359;
        15'h31D1: data = 12'h344;
        15'h31D2: data = 12'h32F;
        15'h31D3: data = 12'h320;
        15'h31D4: data = 12'h30C;
        15'h31D5: data = 12'h2FD;
        15'h31D6: data = 12'h2EF;
        15'h31D7: data = 12'h2DC;
        15'h31D8: data = 12'h2D5;
        15'h31D9: data = 12'h2CF;
        15'h31DA: data = 12'h2C3;
        15'h31DB: data = 12'h2B4;
        15'h31DC: data = 12'h2A7;
        15'h31DD: data = 12'h29E;
        15'h31DE: data = 12'h295;
        15'h31DF: data = 12'h282;
        15'h31E0: data = 12'h27D;
        15'h31E1: data = 12'h26B;
        15'h31E2: data = 12'h262;
        15'h31E3: data = 12'h251;
        15'h31E4: data = 12'h245;
        15'h31E5: data = 12'h230;
        15'h31E6: data = 12'h222;
        15'h31E7: data = 12'h216;
        15'h31E8: data = 12'h20D;
        15'h31E9: data = 12'h207;
        15'h31EA: data = 12'h203;
        15'h31EB: data = 12'h1F6;
        15'h31EC: data = 12'h1F0;
        15'h31ED: data = 12'h1F0;
        15'h31EE: data = 12'h1EA;
        15'h31EF: data = 12'h1E2;
        15'h31F0: data = 12'h1D7;
        15'h31F1: data = 12'h1C9;
        15'h31F2: data = 12'h1C2;
        15'h31F3: data = 12'h1BF;
        15'h31F4: data = 12'h1B4;
        15'h31F5: data = 12'h1A8;
        15'h31F6: data = 12'h19D;
        15'h31F7: data = 12'h191;
        15'h31F8: data = 12'h191;
        15'h31F9: data = 12'h18B;
        15'h31FA: data = 12'h184;
        15'h31FB: data = 12'h183;
        15'h31FC: data = 12'h187;
        15'h31FD: data = 12'h181;
        15'h31FE: data = 12'h185;
        15'h31FF: data = 12'h17E;
        15'h3200: data = 12'h17E;
        15'h3201: data = 12'h177;
        15'h3202: data = 12'h174;
        15'h3203: data = 12'h171;
        15'h3204: data = 12'h165;
        15'h3205: data = 12'h162;
        15'h3206: data = 12'h15D;
        15'h3207: data = 12'h159;
        15'h3208: data = 12'h154;
        15'h3209: data = 12'h155;
        15'h320A: data = 12'h15B;
        15'h320B: data = 12'h15F;
        15'h320C: data = 12'h15F;
        15'h320D: data = 12'h163;
        15'h320E: data = 12'h164;
        15'h320F: data = 12'h170;
        15'h3210: data = 12'h170;
        15'h3211: data = 12'h16F;
        15'h3212: data = 12'h16C;
        15'h3213: data = 12'h167;
        15'h3214: data = 12'h16D;
        15'h3215: data = 12'h16A;
        15'h3216: data = 12'h168;
        15'h3217: data = 12'h16B;
        15'h3218: data = 12'h16A;
        15'h3219: data = 12'h176;
        15'h321A: data = 12'h17C;
        15'h321B: data = 12'h181;
        15'h321C: data = 12'h18D;
        15'h321D: data = 12'h195;
        15'h321E: data = 12'h19C;
        15'h321F: data = 12'h1A6;
        15'h3220: data = 12'h1AB;
        15'h3221: data = 12'h1B4;
        15'h3222: data = 12'h1B2;
        15'h3223: data = 12'h1B9;
        15'h3224: data = 12'h1BA;
        15'h3225: data = 12'h1BD;
        15'h3226: data = 12'h1C7;
        15'h3227: data = 12'h1C8;
        15'h3228: data = 12'h1CF;
        15'h3229: data = 12'h1D5;
        15'h322A: data = 12'h1E1;
        15'h322B: data = 12'h1EE;
        15'h322C: data = 12'h1FB;
        15'h322D: data = 12'h209;
        15'h322E: data = 12'h219;
        15'h322F: data = 12'h21C;
        15'h3230: data = 12'h22C;
        15'h3231: data = 12'h234;
        15'h3232: data = 12'h247;
        15'h3233: data = 12'h24D;
        15'h3234: data = 12'h25C;
        15'h3235: data = 12'h267;
        15'h3236: data = 12'h270;
        15'h3237: data = 12'h272;
        15'h3238: data = 12'h27D;
        15'h3239: data = 12'h28A;
        15'h323A: data = 12'h291;
        15'h323B: data = 12'h29F;
        15'h323C: data = 12'h2B0;
        15'h323D: data = 12'h2C3;
        15'h323E: data = 12'h2CF;
        15'h323F: data = 12'h2DC;
        15'h3240: data = 12'h2EF;
        15'h3241: data = 12'h2FF;
        15'h3242: data = 12'h312;
        15'h3243: data = 12'h326;
        15'h3244: data = 12'h337;
        15'h3245: data = 12'h347;
        15'h3246: data = 12'h355;
        15'h3247: data = 12'h365;
        15'h3248: data = 12'h371;
        15'h3249: data = 12'h380;
        15'h324A: data = 12'h395;
        15'h324B: data = 12'h39A;
        15'h324C: data = 12'h3AC;
        15'h324D: data = 12'h3BB;
        15'h324E: data = 12'h3C6;
        15'h324F: data = 12'h3DB;
        15'h3250: data = 12'h3EE;
        15'h3251: data = 12'h3FB;
        15'h3252: data = 12'h414;
        15'h3253: data = 12'h424;
        15'h3254: data = 12'h43B;
        15'h3255: data = 12'h453;
        15'h3256: data = 12'h467;
        15'h3257: data = 12'h47F;
        15'h3258: data = 12'h48F;
        15'h3259: data = 12'h4A6;
        15'h325A: data = 12'h4B9;
        15'h325B: data = 12'h4CE;
        15'h325C: data = 12'h4E4;
        15'h325D: data = 12'h4F7;
        15'h325E: data = 12'h508;
        15'h325F: data = 12'h51B;
        15'h3260: data = 12'h52C;
        15'h3261: data = 12'h53E;
        15'h3262: data = 12'h553;
        15'h3263: data = 12'h563;
        15'h3264: data = 12'h575;
        15'h3265: data = 12'h58D;
        15'h3266: data = 12'h5A2;
        15'h3267: data = 12'h5B5;
        15'h3268: data = 12'h5CC;
        15'h3269: data = 12'h5E4;
        15'h326A: data = 12'h5FB;
        15'h326B: data = 12'h615;
        15'h326C: data = 12'h62C;
        15'h326D: data = 12'h644;
        15'h326E: data = 12'h65D;
        15'h326F: data = 12'h679;
        15'h3270: data = 12'h68E;
        15'h3271: data = 12'h6A3;
        15'h3272: data = 12'h6B9;
        15'h3273: data = 12'h6D2;
        15'h3274: data = 12'h6E2;
        15'h3275: data = 12'h6F9;
        15'h3276: data = 12'h70C;
        15'h3277: data = 12'h722;
        15'h3278: data = 12'h73A;
        15'h3279: data = 12'h748;
        15'h327A: data = 12'h75F;
        15'h327B: data = 12'h774;
        15'h327C: data = 12'h791;
        15'h327D: data = 12'h7A2;
        15'h327E: data = 12'h7B6;
        15'h327F: data = 12'h7D1;
        15'h3280: data = 12'h7E7;
        15'h3281: data = 12'h800;
        15'h3282: data = 12'h06E;
        15'h3283: data = 12'h085;
        15'h3284: data = 12'h09C;
        15'h3285: data = 12'h0B3;
        15'h3286: data = 12'h0CD;
        15'h3287: data = 12'h0E6;
        15'h3288: data = 12'h100;
        15'h3289: data = 12'h113;
        15'h328A: data = 12'h12A;
        15'h328B: data = 12'h143;
        15'h328C: data = 12'h158;
        15'h328D: data = 12'h16A;
        15'h328E: data = 12'h181;
        15'h328F: data = 12'h19C;
        15'h3290: data = 12'h1B1;
        15'h3291: data = 12'h1C1;
        15'h3292: data = 12'h1D9;
        15'h3293: data = 12'h1EF;
        15'h3294: data = 12'h205;
        15'h3295: data = 12'h218;
        15'h3296: data = 12'h231;
        15'h3297: data = 12'h246;
        15'h3298: data = 12'h25F;
        15'h3299: data = 12'h276;
        15'h329A: data = 12'h28E;
        15'h329B: data = 12'h2A6;
        15'h329C: data = 12'h2BA;
        15'h329D: data = 12'h2D0;
        15'h329E: data = 12'h2ED;
        15'h329F: data = 12'h305;
        15'h32A0: data = 12'h31F;
        15'h32A1: data = 12'h332;
        15'h32A2: data = 12'h34C;
        15'h32A3: data = 12'h367;
        15'h32A4: data = 12'h37C;
        15'h32A5: data = 12'h399;
        15'h32A6: data = 12'h3A8;
        15'h32A7: data = 12'h3C3;
        15'h32A8: data = 12'h3D9;
        15'h32A9: data = 12'h3F0;
        15'h32AA: data = 12'h402;
        15'h32AB: data = 12'h417;
        15'h32AC: data = 12'h42C;
        15'h32AD: data = 12'h442;
        15'h32AE: data = 12'h453;
        15'h32AF: data = 12'h46A;
        15'h32B0: data = 12'h481;
        15'h32B1: data = 12'h496;
        15'h32B2: data = 12'h4AD;
        15'h32B3: data = 12'h4BB;
        15'h32B4: data = 12'h4C9;
        15'h32B5: data = 12'h4DF;
        15'h32B6: data = 12'h4F6;
        15'h32B7: data = 12'h509;
        15'h32B8: data = 12'h517;
        15'h32B9: data = 12'h529;
        15'h32BA: data = 12'h53E;
        15'h32BB: data = 12'h54B;
        15'h32BC: data = 12'h55C;
        15'h32BD: data = 12'h56C;
        15'h32BE: data = 12'h580;
        15'h32BF: data = 12'h590;
        15'h32C0: data = 12'h5A6;
        15'h32C1: data = 12'h5B8;
        15'h32C2: data = 12'h5C4;
        15'h32C3: data = 12'h5D6;
        15'h32C4: data = 12'h5EC;
        15'h32C5: data = 12'h5FA;
        15'h32C6: data = 12'h609;
        15'h32C7: data = 12'h61B;
        15'h32C8: data = 12'h62C;
        15'h32C9: data = 12'h63C;
        15'h32CA: data = 12'h650;
        15'h32CB: data = 12'h65E;
        15'h32CC: data = 12'h66F;
        15'h32CD: data = 12'h67E;
        15'h32CE: data = 12'h691;
        15'h32CF: data = 12'h6A0;
        15'h32D0: data = 12'h6B0;
        15'h32D1: data = 12'h6BF;
        15'h32D2: data = 12'h6D1;
        15'h32D3: data = 12'h6D8;
        15'h32D4: data = 12'h6EA;
        15'h32D5: data = 12'h6FA;
        15'h32D6: data = 12'h709;
        15'h32D7: data = 12'h713;
        15'h32D8: data = 12'h725;
        15'h32D9: data = 12'h731;
        15'h32DA: data = 12'h73B;
        15'h32DB: data = 12'h747;
        15'h32DC: data = 12'h750;
        15'h32DD: data = 12'h75F;
        15'h32DE: data = 12'h767;
        15'h32DF: data = 12'h777;
        15'h32E0: data = 12'h77E;
        15'h32E1: data = 12'h78E;
        15'h32E2: data = 12'h797;
        15'h32E3: data = 12'h79D;
        15'h32E4: data = 12'h7A5;
        15'h32E5: data = 12'h7B1;
        15'h32E6: data = 12'h7B9;
        15'h32E7: data = 12'h7BE;
        15'h32E8: data = 12'h7C8;
        15'h32E9: data = 12'h7CD;
        15'h32EA: data = 12'h7D5;
        15'h32EB: data = 12'h7DD;
        15'h32EC: data = 12'h7E5;
        15'h32ED: data = 12'h7EA;
        15'h32EE: data = 12'h7F2;
        15'h32EF: data = 12'h7FB;
        15'h32F0: data = 12'h7FD;
        15'h32F1: data = 12'h804;
        15'h32F2: data = 12'h807;
        15'h32F3: data = 12'h80D;
        15'h32F4: data = 12'h07B;
        15'h32F5: data = 12'h08B;
        15'h32F6: data = 12'h093;
        15'h32F7: data = 12'h099;
        15'h32F8: data = 12'h09A;
        15'h32F9: data = 12'h0A1;
        15'h32FA: data = 12'h0A0;
        15'h32FB: data = 12'h0A9;
        15'h32FC: data = 12'h0AA;
        15'h32FD: data = 12'h0AD;
        15'h32FE: data = 12'h0B4;
        15'h32FF: data = 12'h0B4;
        15'h3300: data = 12'h0B4;
        15'h3301: data = 12'h0B7;
        15'h3302: data = 12'h0C3;
        15'h3303: data = 12'h0C9;
        15'h3304: data = 12'h0CA;
        15'h3305: data = 12'h0CF;
        15'h3306: data = 12'h0CF;
        15'h3307: data = 12'h0D4;
        15'h3308: data = 12'h0D4;
        15'h3309: data = 12'h0CB;
        15'h330A: data = 12'h0CB;
        15'h330B: data = 12'h0CB;
        15'h330C: data = 12'h0CA;
        15'h330D: data = 12'h0C6;
        15'h330E: data = 12'h0BC;
        15'h330F: data = 12'h0B7;
        15'h3310: data = 12'h0AE;
        15'h3311: data = 12'h0AD;
        15'h3312: data = 12'h0A4;
        15'h3313: data = 12'h0A7;
        15'h3314: data = 12'h0A7;
        15'h3315: data = 12'h0AE;
        15'h3316: data = 12'h0AC;
        15'h3317: data = 12'h0A1;
        15'h3318: data = 12'h0A7;
        15'h3319: data = 12'h099;
        15'h331A: data = 12'h092;
        15'h331B: data = 12'h083;
        15'h331C: data = 12'h077;
        15'h331D: data = 12'h074;
        15'h331E: data = 12'h06D;
        15'h331F: data = 12'h069;
        15'h3320: data = 12'h065;
        15'h3321: data = 12'h063;
        15'h3322: data = 12'h060;
        15'h3323: data = 12'h055;
        15'h3324: data = 12'h046;
        15'h3325: data = 12'h7C4;
        15'h3326: data = 12'h7B3;
        15'h3327: data = 12'h7A7;
        15'h3328: data = 12'h79B;
        15'h3329: data = 12'h794;
        15'h332A: data = 12'h78E;
        15'h332B: data = 12'h788;
        15'h332C: data = 12'h77D;
        15'h332D: data = 12'h76F;
        15'h332E: data = 12'h75E;
        15'h332F: data = 12'h747;
        15'h3330: data = 12'h73B;
        15'h3331: data = 12'h72D;
        15'h3332: data = 12'h723;
        15'h3333: data = 12'h718;
        15'h3334: data = 12'h70E;
        15'h3335: data = 12'h709;
        15'h3336: data = 12'h6FC;
        15'h3337: data = 12'h6EE;
        15'h3338: data = 12'h6DE;
        15'h3339: data = 12'h6D0;
        15'h333A: data = 12'h6B7;
        15'h333B: data = 12'h6A4;
        15'h333C: data = 12'h696;
        15'h333D: data = 12'h686;
        15'h333E: data = 12'h67A;
        15'h333F: data = 12'h66D;
        15'h3340: data = 12'h661;
        15'h3341: data = 12'h653;
        15'h3342: data = 12'h646;
        15'h3343: data = 12'h635;
        15'h3344: data = 12'h62F;
        15'h3345: data = 12'h614;
        15'h3346: data = 12'h605;
        15'h3347: data = 12'h5EB;
        15'h3348: data = 12'h5D0;
        15'h3349: data = 12'h5C0;
        15'h334A: data = 12'h5B0;
        15'h334B: data = 12'h59F;
        15'h334C: data = 12'h58D;
        15'h334D: data = 12'h57A;
        15'h334E: data = 12'h568;
        15'h334F: data = 12'h55D;
        15'h3350: data = 12'h550;
        15'h3351: data = 12'h53F;
        15'h3352: data = 12'h52B;
        15'h3353: data = 12'h518;
        15'h3354: data = 12'h507;
        15'h3355: data = 12'h4F7;
        15'h3356: data = 12'h4DB;
        15'h3357: data = 12'h4C9;
        15'h3358: data = 12'h4B6;
        15'h3359: data = 12'h49B;
        15'h335A: data = 12'h486;
        15'h335B: data = 12'h46D;
        15'h335C: data = 12'h459;
        15'h335D: data = 12'h441;
        15'h335E: data = 12'h429;
        15'h335F: data = 12'h416;
        15'h3360: data = 12'h3FE;
        15'h3361: data = 12'h3E8;
        15'h3362: data = 12'h3D3;
        15'h3363: data = 12'h3C1;
        15'h3364: data = 12'h3AE;
        15'h3365: data = 12'h38F;
        15'h3366: data = 12'h37C;
        15'h3367: data = 12'h365;
        15'h3368: data = 12'h352;
        15'h3369: data = 12'h33D;
        15'h336A: data = 12'h327;
        15'h336B: data = 12'h313;
        15'h336C: data = 12'h2F9;
        15'h336D: data = 12'h2E2;
        15'h336E: data = 12'h2D2;
        15'h336F: data = 12'h2BA;
        15'h3370: data = 12'h2A7;
        15'h3371: data = 12'h289;
        15'h3372: data = 12'h27C;
        15'h3373: data = 12'h261;
        15'h3374: data = 12'h246;
        15'h3375: data = 12'h231;
        15'h3376: data = 12'h218;
        15'h3377: data = 12'h203;
        15'h3378: data = 12'h1F1;
        15'h3379: data = 12'h1D4;
        15'h337A: data = 12'h1BE;
        15'h337B: data = 12'h1A7;
        15'h337C: data = 12'h195;
        15'h337D: data = 12'h179;
        15'h337E: data = 12'h166;
        15'h337F: data = 12'h14C;
        15'h3380: data = 12'h136;
        15'h3381: data = 12'h11D;
        15'h3382: data = 12'h10A;
        15'h3383: data = 12'h0F3;
        15'h3384: data = 12'h0DA;
        15'h3385: data = 12'h0BD;
        15'h3386: data = 12'h0A7;
        15'h3387: data = 12'h090;
        15'h3388: data = 12'h07C;
        15'h3389: data = 12'h065;
        15'h338A: data = 12'h04D;
        15'h338B: data = 12'h7E4;
        15'h338C: data = 12'h7CE;
        15'h338D: data = 12'h7B9;
        15'h338E: data = 12'h7A4;
        15'h338F: data = 12'h78C;
        15'h3390: data = 12'h778;
        15'h3391: data = 12'h75C;
        15'h3392: data = 12'h74C;
        15'h3393: data = 12'h734;
        15'h3394: data = 12'h71E;
        15'h3395: data = 12'h70A;
        15'h3396: data = 12'h6ED;
        15'h3397: data = 12'h6D9;
        15'h3398: data = 12'h6C6;
        15'h3399: data = 12'h6AF;
        15'h339A: data = 12'h695;
        15'h339B: data = 12'h682;
        15'h339C: data = 12'h669;
        15'h339D: data = 12'h655;
        15'h339E: data = 12'h63B;
        15'h339F: data = 12'h628;
        15'h33A0: data = 12'h615;
        15'h33A1: data = 12'h5FA;
        15'h33A2: data = 12'h5E6;
        15'h33A3: data = 12'h5D0;
        15'h33A4: data = 12'h5BD;
        15'h33A5: data = 12'h5A0;
        15'h33A6: data = 12'h588;
        15'h33A7: data = 12'h573;
        15'h33A8: data = 12'h561;
        15'h33A9: data = 12'h54C;
        15'h33AA: data = 12'h536;
        15'h33AB: data = 12'h51C;
        15'h33AC: data = 12'h508;
        15'h33AD: data = 12'h4F5;
        15'h33AE: data = 12'h4DE;
        15'h33AF: data = 12'h4CA;
        15'h33B0: data = 12'h4B6;
        15'h33B1: data = 12'h4A3;
        15'h33B2: data = 12'h48D;
        15'h33B3: data = 12'h47E;
        15'h33B4: data = 12'h466;
        15'h33B5: data = 12'h453;
        15'h33B6: data = 12'h447;
        15'h33B7: data = 12'h435;
        15'h33B8: data = 12'h423;
        15'h33B9: data = 12'h416;
        15'h33BA: data = 12'h401;
        15'h33BB: data = 12'h3F4;
        15'h33BC: data = 12'h3E7;
        15'h33BD: data = 12'h3D2;
        15'h33BE: data = 12'h3C3;
        15'h33BF: data = 12'h3B3;
        15'h33C0: data = 12'h39C;
        15'h33C1: data = 12'h392;
        15'h33C2: data = 12'h378;
        15'h33C3: data = 12'h368;
        15'h33C4: data = 12'h357;
        15'h33C5: data = 12'h346;
        15'h33C6: data = 12'h331;
        15'h33C7: data = 12'h31F;
        15'h33C8: data = 12'h30E;
        15'h33C9: data = 12'h2FD;
        15'h33CA: data = 12'h2F0;
        15'h33CB: data = 12'h2E0;
        15'h33CC: data = 12'h2D3;
        15'h33CD: data = 12'h2CE;
        15'h33CE: data = 12'h2C3;
        15'h33CF: data = 12'h2B5;
        15'h33D0: data = 12'h2A9;
        15'h33D1: data = 12'h29E;
        15'h33D2: data = 12'h293;
        15'h33D3: data = 12'h287;
        15'h33D4: data = 12'h27D;
        15'h33D5: data = 12'h26E;
        15'h33D6: data = 12'h263;
        15'h33D7: data = 12'h251;
        15'h33D8: data = 12'h245;
        15'h33D9: data = 12'h235;
        15'h33DA: data = 12'h222;
        15'h33DB: data = 12'h215;
        15'h33DC: data = 12'h20E;
        15'h33DD: data = 12'h206;
        15'h33DE: data = 12'h201;
        15'h33DF: data = 12'h1F1;
        15'h33E0: data = 12'h1F1;
        15'h33E1: data = 12'h1EF;
        15'h33E2: data = 12'h1E9;
        15'h33E3: data = 12'h1E2;
        15'h33E4: data = 12'h1D4;
        15'h33E5: data = 12'h1CC;
        15'h33E6: data = 12'h1C2;
        15'h33E7: data = 12'h1BE;
        15'h33E8: data = 12'h1B7;
        15'h33E9: data = 12'h1A7;
        15'h33EA: data = 12'h19D;
        15'h33EB: data = 12'h191;
        15'h33EC: data = 12'h191;
        15'h33ED: data = 12'h189;
        15'h33EE: data = 12'h185;
        15'h33EF: data = 12'h185;
        15'h33F0: data = 12'h186;
        15'h33F1: data = 12'h182;
        15'h33F2: data = 12'h185;
        15'h33F3: data = 12'h17F;
        15'h33F4: data = 12'h180;
        15'h33F5: data = 12'h175;
        15'h33F6: data = 12'h174;
        15'h33F7: data = 12'h173;
        15'h33F8: data = 12'h167;
        15'h33F9: data = 12'h162;
        15'h33FA: data = 12'h15C;
        15'h33FB: data = 12'h15E;
        15'h33FC: data = 12'h155;
        15'h33FD: data = 12'h156;
        15'h33FE: data = 12'h159;
        15'h33FF: data = 12'h15B;
        15'h3400: data = 12'h15F;
        15'h3401: data = 12'h164;
        15'h3402: data = 12'h167;
        15'h3403: data = 12'h171;
        15'h3404: data = 12'h16F;
        15'h3405: data = 12'h16F;
        15'h3406: data = 12'h16D;
        15'h3407: data = 12'h16B;
        15'h3408: data = 12'h16F;
        15'h3409: data = 12'h16B;
        15'h340A: data = 12'h16C;
        15'h340B: data = 12'h16D;
        15'h340C: data = 12'h16A;
        15'h340D: data = 12'h176;
        15'h340E: data = 12'h17F;
        15'h340F: data = 12'h183;
        15'h3410: data = 12'h18B;
        15'h3411: data = 12'h18F;
        15'h3412: data = 12'h19B;
        15'h3413: data = 12'h1A2;
        15'h3414: data = 12'h1AE;
        15'h3415: data = 12'h1B3;
        15'h3416: data = 12'h1B4;
        15'h3417: data = 12'h1BB;
        15'h3418: data = 12'h1C1;
        15'h3419: data = 12'h1C2;
        15'h341A: data = 12'h1C2;
        15'h341B: data = 12'h1CB;
        15'h341C: data = 12'h1D1;
        15'h341D: data = 12'h1D7;
        15'h341E: data = 12'h1E1;
        15'h341F: data = 12'h1F1;
        15'h3420: data = 12'h1FA;
        15'h3421: data = 12'h203;
        15'h3422: data = 12'h218;
        15'h3423: data = 12'h21D;
        15'h3424: data = 12'h230;
        15'h3425: data = 12'h239;
        15'h3426: data = 12'h247;
        15'h3427: data = 12'h24F;
        15'h3428: data = 12'h25C;
        15'h3429: data = 12'h265;
        15'h342A: data = 12'h26F;
        15'h342B: data = 12'h273;
        15'h342C: data = 12'h280;
        15'h342D: data = 12'h28A;
        15'h342E: data = 12'h291;
        15'h342F: data = 12'h29F;
        15'h3430: data = 12'h2B2;
        15'h3431: data = 12'h2BF;
        15'h3432: data = 12'h2D1;
        15'h3433: data = 12'h2DD;
        15'h3434: data = 12'h2EF;
        15'h3435: data = 12'h2FF;
        15'h3436: data = 12'h310;
        15'h3437: data = 12'h326;
        15'h3438: data = 12'h338;
        15'h3439: data = 12'h345;
        15'h343A: data = 12'h357;
        15'h343B: data = 12'h363;
        15'h343C: data = 12'h373;
        15'h343D: data = 12'h380;
        15'h343E: data = 12'h396;
        15'h343F: data = 12'h39C;
        15'h3440: data = 12'h3B0;
        15'h3441: data = 12'h3BB;
        15'h3442: data = 12'h3CB;
        15'h3443: data = 12'h3DD;
        15'h3444: data = 12'h3EE;
        15'h3445: data = 12'h3FD;
        15'h3446: data = 12'h412;
        15'h3447: data = 12'h428;
        15'h3448: data = 12'h43E;
        15'h3449: data = 12'h453;
        15'h344A: data = 12'h466;
        15'h344B: data = 12'h47F;
        15'h344C: data = 12'h494;
        15'h344D: data = 12'h4AC;
        15'h344E: data = 12'h4B8;
        15'h344F: data = 12'h4D1;
        15'h3450: data = 12'h4E4;
        15'h3451: data = 12'h4F9;
        15'h3452: data = 12'h511;
        15'h3453: data = 12'h51F;
        15'h3454: data = 12'h52F;
        15'h3455: data = 12'h544;
        15'h3456: data = 12'h556;
        15'h3457: data = 12'h568;
        15'h3458: data = 12'h577;
        15'h3459: data = 12'h58B;
        15'h345A: data = 12'h5A3;
        15'h345B: data = 12'h5B4;
        15'h345C: data = 12'h5CB;
        15'h345D: data = 12'h5E3;
        15'h345E: data = 12'h5F6;
        15'h345F: data = 12'h614;
        15'h3460: data = 12'h62D;
        15'h3461: data = 12'h646;
        15'h3462: data = 12'h662;
        15'h3463: data = 12'h676;
        15'h3464: data = 12'h692;
        15'h3465: data = 12'h6A2;
        15'h3466: data = 12'h6BA;
        15'h3467: data = 12'h6D4;
        15'h3468: data = 12'h6E3;
        15'h3469: data = 12'h6F9;
        15'h346A: data = 12'h70F;
        15'h346B: data = 12'h721;
        15'h346C: data = 12'h739;
        15'h346D: data = 12'h749;
        15'h346E: data = 12'h761;
        15'h346F: data = 12'h777;
        15'h3470: data = 12'h790;
        15'h3471: data = 12'h79E;
        15'h3472: data = 12'h7B8;
        15'h3473: data = 12'h7D3;
        15'h3474: data = 12'h7E8;
        15'h3475: data = 12'h800;
        15'h3476: data = 12'h071;
        15'h3477: data = 12'h085;
        15'h3478: data = 12'h09F;
        15'h3479: data = 12'h0B5;
        15'h347A: data = 12'h0D3;
        15'h347B: data = 12'h0E9;
        15'h347C: data = 12'h103;
        15'h347D: data = 12'h117;
        15'h347E: data = 12'h12C;
        15'h347F: data = 12'h145;
        15'h3480: data = 12'h158;
        15'h3481: data = 12'h170;
        15'h3482: data = 12'h185;
        15'h3483: data = 12'h19F;
        15'h3484: data = 12'h1B5;
        15'h3485: data = 12'h1C2;
        15'h3486: data = 12'h1DE;
        15'h3487: data = 12'h1F4;
        15'h3488: data = 12'h209;
        15'h3489: data = 12'h21A;
        15'h348A: data = 12'h234;
        15'h348B: data = 12'h248;
        15'h348C: data = 12'h262;
        15'h348D: data = 12'h273;
        15'h348E: data = 12'h28F;
        15'h348F: data = 12'h2A3;
        15'h3490: data = 12'h2BD;
        15'h3491: data = 12'h2D2;
        15'h3492: data = 12'h2EA;
        15'h3493: data = 12'h308;
        15'h3494: data = 12'h31F;
        15'h3495: data = 12'h334;
        15'h3496: data = 12'h347;
        15'h3497: data = 12'h366;
        15'h3498: data = 12'h379;
        15'h3499: data = 12'h395;
        15'h349A: data = 12'h3A7;
        15'h349B: data = 12'h3C0;
        15'h349C: data = 12'h3DA;
        15'h349D: data = 12'h3ED;
        15'h349E: data = 12'h401;
        15'h349F: data = 12'h418;
        15'h34A0: data = 12'h42E;
        15'h34A1: data = 12'h445;
        15'h34A2: data = 12'h454;
        15'h34A3: data = 12'h469;
        15'h34A4: data = 12'h481;
        15'h34A5: data = 12'h497;
        15'h34A6: data = 12'h4AC;
        15'h34A7: data = 12'h4B8;
        15'h34A8: data = 12'h4CA;
        15'h34A9: data = 12'h4DF;
        15'h34AA: data = 12'h4F5;
        15'h34AB: data = 12'h50A;
        15'h34AC: data = 12'h515;
        15'h34AD: data = 12'h52A;
        15'h34AE: data = 12'h53C;
        15'h34AF: data = 12'h54C;
        15'h34B0: data = 12'h55D;
        15'h34B1: data = 12'h56E;
        15'h34B2: data = 12'h582;
        15'h34B3: data = 12'h591;
        15'h34B4: data = 12'h5A5;
        15'h34B5: data = 12'h5B7;
        15'h34B6: data = 12'h5C4;
        15'h34B7: data = 12'h5D6;
        15'h34B8: data = 12'h5E9;
        15'h34B9: data = 12'h5FC;
        15'h34BA: data = 12'h60C;
        15'h34BB: data = 12'h618;
        15'h34BC: data = 12'h62A;
        15'h34BD: data = 12'h63A;
        15'h34BE: data = 12'h64F;
        15'h34BF: data = 12'h65D;
        15'h34C0: data = 12'h670;
        15'h34C1: data = 12'h680;
        15'h34C2: data = 12'h691;
        15'h34C3: data = 12'h6A0;
        15'h34C4: data = 12'h6AE;
        15'h34C5: data = 12'h6C1;
        15'h34C6: data = 12'h6CE;
        15'h34C7: data = 12'h6D8;
        15'h34C8: data = 12'h6EB;
        15'h34C9: data = 12'h6F8;
        15'h34CA: data = 12'h705;
        15'h34CB: data = 12'h712;
        15'h34CC: data = 12'h723;
        15'h34CD: data = 12'h732;
        15'h34CE: data = 12'h736;
        15'h34CF: data = 12'h743;
        15'h34D0: data = 12'h750;
        15'h34D1: data = 12'h75F;
        15'h34D2: data = 12'h767;
        15'h34D3: data = 12'h778;
        15'h34D4: data = 12'h77D;
        15'h34D5: data = 12'h78D;
        15'h34D6: data = 12'h794;
        15'h34D7: data = 12'h79F;
        15'h34D8: data = 12'h7A4;
        15'h34D9: data = 12'h7AF;
        15'h34DA: data = 12'h7BA;
        15'h34DB: data = 12'h7BD;
        15'h34DC: data = 12'h7C8;
        15'h34DD: data = 12'h7CE;
        15'h34DE: data = 12'h7D4;
        15'h34DF: data = 12'h7DE;
        15'h34E0: data = 12'h7EA;
        15'h34E1: data = 12'h7E8;
        15'h34E2: data = 12'h7F4;
        15'h34E3: data = 12'h7FB;
        15'h34E4: data = 12'h802;
        15'h34E5: data = 12'h806;
        15'h34E6: data = 12'h805;
        15'h34E7: data = 12'h80B;
        15'h34E8: data = 12'h812;
        15'h34E9: data = 12'h08F;
        15'h34EA: data = 12'h095;
        15'h34EB: data = 12'h09B;
        15'h34EC: data = 12'h09D;
        15'h34ED: data = 12'h0A5;
        15'h34EE: data = 12'h0A3;
        15'h34EF: data = 12'h0AC;
        15'h34F0: data = 12'h0AD;
        15'h34F1: data = 12'h0AA;
        15'h34F2: data = 12'h0B5;
        15'h34F3: data = 12'h0B5;
        15'h34F4: data = 12'h0B6;
        15'h34F5: data = 12'h0B9;
        15'h34F6: data = 12'h0C2;
        15'h34F7: data = 12'h0C3;
        15'h34F8: data = 12'h0C5;
        15'h34F9: data = 12'h0CA;
        15'h34FA: data = 12'h0CB;
        15'h34FB: data = 12'h0D0;
        15'h34FC: data = 12'h0D6;
        15'h34FD: data = 12'h0CE;
        15'h34FE: data = 12'h0D0;
        15'h34FF: data = 12'h0CE;
        15'h3500: data = 12'h0CB;
        15'h3501: data = 12'h0C8;
        15'h3502: data = 12'h0BF;
        15'h3503: data = 12'h0BC;
        15'h3504: data = 12'h0B1;
        15'h3505: data = 12'h0AD;
        15'h3506: data = 12'h0A3;
        15'h3507: data = 12'h0A5;
        15'h3508: data = 12'h0A0;
        15'h3509: data = 12'h0A9;
        15'h350A: data = 12'h0A9;
        15'h350B: data = 12'h0A5;
        15'h350C: data = 12'h0A7;
        15'h350D: data = 12'h09D;
        15'h350E: data = 12'h090;
        15'h350F: data = 12'h085;
        15'h3510: data = 12'h078;
        15'h3511: data = 12'h075;
        15'h3512: data = 12'h06B;
        15'h3513: data = 12'h065;
        15'h3514: data = 12'h064;
        15'h3515: data = 12'h065;
        15'h3516: data = 12'h061;
        15'h3517: data = 12'h055;
        15'h3518: data = 12'h049;
        15'h3519: data = 12'h443;
        15'h351A: data = 12'h7B9;
        15'h351B: data = 12'h7AB;
        15'h351C: data = 12'h79E;
        15'h351D: data = 12'h790;
        15'h351E: data = 12'h78C;
        15'h351F: data = 12'h788;
        15'h3520: data = 12'h77C;
        15'h3521: data = 12'h770;
        15'h3522: data = 12'h761;
        15'h3523: data = 12'h74C;
        15'h3524: data = 12'h73B;
        15'h3525: data = 12'h72E;
        15'h3526: data = 12'h722;
        15'h3527: data = 12'h714;
        15'h3528: data = 12'h70D;
        15'h3529: data = 12'h708;
        15'h352A: data = 12'h6FA;
        15'h352B: data = 12'h6EA;
        15'h352C: data = 12'h6DF;
        15'h352D: data = 12'h6CE;
        15'h352E: data = 12'h6BA;
        15'h352F: data = 12'h6AA;
        15'h3530: data = 12'h693;
        15'h3531: data = 12'h685;
        15'h3532: data = 12'h678;
        15'h3533: data = 12'h66F;
        15'h3534: data = 12'h661;
        15'h3535: data = 12'h658;
        15'h3536: data = 12'h649;
        15'h3537: data = 12'h635;
        15'h3538: data = 12'h62B;
        15'h3539: data = 12'h614;
        15'h353A: data = 12'h605;
        15'h353B: data = 12'h5F0;
        15'h353C: data = 12'h5D1;
        15'h353D: data = 12'h5C2;
        15'h353E: data = 12'h5B4;
        15'h353F: data = 12'h59E;
        15'h3540: data = 12'h58E;
        15'h3541: data = 12'h57B;
        15'h3542: data = 12'h56D;
        15'h3543: data = 12'h55F;
        15'h3544: data = 12'h554;
        15'h3545: data = 12'h542;
        15'h3546: data = 12'h529;
        15'h3547: data = 12'h51A;
        15'h3548: data = 12'h505;
        15'h3549: data = 12'h4F7;
        15'h354A: data = 12'h4DE;
        15'h354B: data = 12'h4C8;
        15'h354C: data = 12'h4B9;
        15'h354D: data = 12'h49D;
        15'h354E: data = 12'h483;
        15'h354F: data = 12'h46C;
        15'h3550: data = 12'h455;
        15'h3551: data = 12'h442;
        15'h3552: data = 12'h42B;
        15'h3553: data = 12'h415;
        15'h3554: data = 12'h3FC;
        15'h3555: data = 12'h3E5;
        15'h3556: data = 12'h3D2;
        15'h3557: data = 12'h3BE;
        15'h3558: data = 12'h3AA;
        15'h3559: data = 12'h391;
        15'h355A: data = 12'h37F;
        15'h355B: data = 12'h36A;
        15'h355C: data = 12'h354;
        15'h355D: data = 12'h33A;
        15'h355E: data = 12'h327;
        15'h355F: data = 12'h314;
        15'h3560: data = 12'h2FC;
        15'h3561: data = 12'h2E9;
        15'h3562: data = 12'h2D5;
        15'h3563: data = 12'h2BF;
        15'h3564: data = 12'h2A3;
        15'h3565: data = 12'h28D;
        15'h3566: data = 12'h27F;
        15'h3567: data = 12'h262;
        15'h3568: data = 12'h24A;
        15'h3569: data = 12'h234;
        15'h356A: data = 12'h21E;
        15'h356B: data = 12'h203;
        15'h356C: data = 12'h1F2;
        15'h356D: data = 12'h1D5;
        15'h356E: data = 12'h1C1;
        15'h356F: data = 12'h1AC;
        15'h3570: data = 12'h195;
        15'h3571: data = 12'h17C;
        15'h3572: data = 12'h167;
        15'h3573: data = 12'h14E;
        15'h3574: data = 12'h138;
        15'h3575: data = 12'h11B;
        15'h3576: data = 12'h109;
        15'h3577: data = 12'h0F6;
        15'h3578: data = 12'h0DB;
        15'h3579: data = 12'h0BE;
        15'h357A: data = 12'h0A7;
        15'h357B: data = 12'h092;
        15'h357C: data = 12'h07E;
        15'h357D: data = 12'h063;
        15'h357E: data = 12'h050;
        15'h357F: data = 12'h7E2;
        15'h3580: data = 12'h7CE;
        15'h3581: data = 12'h7BD;
        15'h3582: data = 12'h7A4;
        15'h3583: data = 12'h78F;
        15'h3584: data = 12'h778;
        15'h3585: data = 12'h75C;
        15'h3586: data = 12'h74B;
        15'h3587: data = 12'h736;
        15'h3588: data = 12'h720;
        15'h3589: data = 12'h70A;
        15'h358A: data = 12'h6EC;
        15'h358B: data = 12'h6DB;
        15'h358C: data = 12'h6C8;
        15'h358D: data = 12'h6B2;
        15'h358E: data = 12'h695;
        15'h358F: data = 12'h67E;
        15'h3590: data = 12'h669;
        15'h3591: data = 12'h652;
        15'h3592: data = 12'h63D;
        15'h3593: data = 12'h62D;
        15'h3594: data = 12'h617;
        15'h3595: data = 12'h5FB;
        15'h3596: data = 12'h5E5;
        15'h3597: data = 12'h5CF;
        15'h3598: data = 12'h5BA;
        15'h3599: data = 12'h59E;
        15'h359A: data = 12'h589;
        15'h359B: data = 12'h572;
        15'h359C: data = 12'h565;
        15'h359D: data = 12'h54A;
        15'h359E: data = 12'h533;
        15'h359F: data = 12'h520;
        15'h35A0: data = 12'h508;
        15'h35A1: data = 12'h4F4;
        15'h35A2: data = 12'h4DB;
        15'h35A3: data = 12'h4C7;
        15'h35A4: data = 12'h4B5;
        15'h35A5: data = 12'h4A2;
        15'h35A6: data = 12'h490;
        15'h35A7: data = 12'h47D;
        15'h35A8: data = 12'h466;
        15'h35A9: data = 12'h456;
        15'h35AA: data = 12'h449;
        15'h35AB: data = 12'h436;
        15'h35AC: data = 12'h423;
        15'h35AD: data = 12'h414;
        15'h35AE: data = 12'h403;
        15'h35AF: data = 12'h3F5;
        15'h35B0: data = 12'h3E6;
        15'h35B1: data = 12'h3D3;
        15'h35B2: data = 12'h3C5;
        15'h35B3: data = 12'h3B0;
        15'h35B4: data = 12'h39A;
        15'h35B5: data = 12'h392;
        15'h35B6: data = 12'h378;
        15'h35B7: data = 12'h369;
        15'h35B8: data = 12'h356;
        15'h35B9: data = 12'h346;
        15'h35BA: data = 12'h333;
        15'h35BB: data = 12'h31F;
        15'h35BC: data = 12'h30D;
        15'h35BD: data = 12'h2FA;
        15'h35BE: data = 12'h2F1;
        15'h35BF: data = 12'h2DF;
        15'h35C0: data = 12'h2D3;
        15'h35C1: data = 12'h2CE;
        15'h35C2: data = 12'h2C1;
        15'h35C3: data = 12'h2B6;
        15'h35C4: data = 12'h2AA;
        15'h35C5: data = 12'h29E;
        15'h35C6: data = 12'h297;
        15'h35C7: data = 12'h285;
        15'h35C8: data = 12'h27D;
        15'h35C9: data = 12'h26C;
        15'h35CA: data = 12'h264;
        15'h35CB: data = 12'h251;
        15'h35CC: data = 12'h241;
        15'h35CD: data = 12'h232;
        15'h35CE: data = 12'h222;
        15'h35CF: data = 12'h213;
        15'h35D0: data = 12'h20F;
        15'h35D1: data = 12'h207;
        15'h35D2: data = 12'h1FF;
        15'h35D3: data = 12'h1F4;
        15'h35D4: data = 12'h1F1;
        15'h35D5: data = 12'h1EE;
        15'h35D6: data = 12'h1EA;
        15'h35D7: data = 12'h1E3;
        15'h35D8: data = 12'h1D4;
        15'h35D9: data = 12'h1C9;
        15'h35DA: data = 12'h1C2;
        15'h35DB: data = 12'h1C0;
        15'h35DC: data = 12'h1B5;
        15'h35DD: data = 12'h1A5;
        15'h35DE: data = 12'h19D;
        15'h35DF: data = 12'h18E;
        15'h35E0: data = 12'h191;
        15'h35E1: data = 12'h18A;
        15'h35E2: data = 12'h188;
        15'h35E3: data = 12'h185;
        15'h35E4: data = 12'h186;
        15'h35E5: data = 12'h186;
        15'h35E6: data = 12'h186;
        15'h35E7: data = 12'h17E;
        15'h35E8: data = 12'h17D;
        15'h35E9: data = 12'h174;
        15'h35EA: data = 12'h171;
        15'h35EB: data = 12'h171;
        15'h35EC: data = 12'h165;
        15'h35ED: data = 12'h161;
        15'h35EE: data = 12'h160;
        15'h35EF: data = 12'h15D;
        15'h35F0: data = 12'h158;
        15'h35F1: data = 12'h156;
        15'h35F2: data = 12'h158;
        15'h35F3: data = 12'h15B;
        15'h35F4: data = 12'h163;
        15'h35F5: data = 12'h163;
        15'h35F6: data = 12'h168;
        15'h35F7: data = 12'h170;
        15'h35F8: data = 12'h16F;
        15'h35F9: data = 12'h16E;
        15'h35FA: data = 12'h16C;
        15'h35FB: data = 12'h16B;
        15'h35FC: data = 12'h16E;
        15'h35FD: data = 12'h16C;
        15'h35FE: data = 12'h16C;
        15'h35FF: data = 12'h16B;
        15'h3600: data = 12'h16A;
        15'h3601: data = 12'h172;
        15'h3602: data = 12'h17D;
        15'h3603: data = 12'h17F;
        15'h3604: data = 12'h188;
        15'h3605: data = 12'h192;
        15'h3606: data = 12'h19B;
        15'h3607: data = 12'h1A6;
        15'h3608: data = 12'h1AE;
        15'h3609: data = 12'h1B4;
        15'h360A: data = 12'h1B4;
        15'h360B: data = 12'h1B9;
        15'h360C: data = 12'h1BD;
        15'h360D: data = 12'h1C3;
        15'h360E: data = 12'h1C5;
        15'h360F: data = 12'h1C8;
        15'h3610: data = 12'h1D3;
        15'h3611: data = 12'h1D8;
        15'h3612: data = 12'h1E3;
        15'h3613: data = 12'h1EE;
        15'h3614: data = 12'h1F9;
        15'h3615: data = 12'h206;
        15'h3616: data = 12'h219;
        15'h3617: data = 12'h21D;
        15'h3618: data = 12'h22D;
        15'h3619: data = 12'h238;
        15'h361A: data = 12'h248;
        15'h361B: data = 12'h24F;
        15'h361C: data = 12'h25C;
        15'h361D: data = 12'h265;
        15'h361E: data = 12'h272;
        15'h361F: data = 12'h273;
        15'h3620: data = 12'h280;
        15'h3621: data = 12'h28C;
        15'h3622: data = 12'h294;
        15'h3623: data = 12'h29F;
        15'h3624: data = 12'h2B0;
        15'h3625: data = 12'h2C2;
        15'h3626: data = 12'h2D2;
        15'h3627: data = 12'h2DA;
        15'h3628: data = 12'h2F0;
        15'h3629: data = 12'h301;
        15'h362A: data = 12'h312;
        15'h362B: data = 12'h325;
        15'h362C: data = 12'h337;
        15'h362D: data = 12'h345;
        15'h362E: data = 12'h358;
        15'h362F: data = 12'h364;
        15'h3630: data = 12'h378;
        15'h3631: data = 12'h37F;
        15'h3632: data = 12'h398;
        15'h3633: data = 12'h39D;
        15'h3634: data = 12'h3B1;
        15'h3635: data = 12'h3BB;
        15'h3636: data = 12'h3C8;
        15'h3637: data = 12'h3DD;
        15'h3638: data = 12'h3EC;
        15'h3639: data = 12'h3FB;
        15'h363A: data = 12'h416;
        15'h363B: data = 12'h429;
        15'h363C: data = 12'h43F;
        15'h363D: data = 12'h456;
        15'h363E: data = 12'h466;
        15'h363F: data = 12'h47D;
        15'h3640: data = 12'h492;
        15'h3641: data = 12'h4A8;
        15'h3642: data = 12'h4BC;
        15'h3643: data = 12'h4D1;
        15'h3644: data = 12'h4E5;
        15'h3645: data = 12'h4F7;
        15'h3646: data = 12'h50B;
        15'h3647: data = 12'h520;
        15'h3648: data = 12'h52D;
        15'h3649: data = 12'h542;
        15'h364A: data = 12'h556;
        15'h364B: data = 12'h567;
        15'h364C: data = 12'h574;
        15'h364D: data = 12'h58E;
        15'h364E: data = 12'h5A2;
        15'h364F: data = 12'h5B6;
        15'h3650: data = 12'h5CA;
        15'h3651: data = 12'h5E2;
        15'h3652: data = 12'h5FA;
        15'h3653: data = 12'h614;
        15'h3654: data = 12'h62B;
        15'h3655: data = 12'h645;
        15'h3656: data = 12'h65D;
        15'h3657: data = 12'h676;
        15'h3658: data = 12'h692;
        15'h3659: data = 12'h6A2;
        15'h365A: data = 12'h6B7;
        15'h365B: data = 12'h6D1;
        15'h365C: data = 12'h6E5;
        15'h365D: data = 12'h6FA;
        15'h365E: data = 12'h70D;
        15'h365F: data = 12'h722;
        15'h3660: data = 12'h73C;
        15'h3661: data = 12'h748;
        15'h3662: data = 12'h75F;
        15'h3663: data = 12'h776;
        15'h3664: data = 12'h78E;
        15'h3665: data = 12'h7A0;
        15'h3666: data = 12'h7B6;
        15'h3667: data = 12'h7D1;
        15'h3668: data = 12'h7E6;
        15'h3669: data = 12'h7FD;
        15'h366A: data = 12'h06E;
        15'h366B: data = 12'h083;
        15'h366C: data = 12'h09C;
        15'h366D: data = 12'h0B0;
        15'h366E: data = 12'h0D0;
        15'h366F: data = 12'h0E9;
        15'h3670: data = 12'h0FF;
        15'h3671: data = 12'h116;
        15'h3672: data = 12'h12C;
        15'h3673: data = 12'h146;
        15'h3674: data = 12'h157;
        15'h3675: data = 12'h171;
        15'h3676: data = 12'h185;
        15'h3677: data = 12'h19F;
        15'h3678: data = 12'h1B5;
        15'h3679: data = 12'h1C1;
        15'h367A: data = 12'h1DE;
        15'h367B: data = 12'h1F3;
        15'h367C: data = 12'h209;
        15'h367D: data = 12'h21C;
        15'h367E: data = 12'h231;
        15'h367F: data = 12'h24A;
        15'h3680: data = 12'h25E;
        15'h3681: data = 12'h274;
        15'h3682: data = 12'h28C;
        15'h3683: data = 12'h2A5;
        15'h3684: data = 12'h2BE;
        15'h3685: data = 12'h2D4;
        15'h3686: data = 12'h2EE;
        15'h3687: data = 12'h305;
        15'h3688: data = 12'h31F;
        15'h3689: data = 12'h332;
        15'h368A: data = 12'h348;
        15'h368B: data = 12'h364;
        15'h368C: data = 12'h378;
        15'h368D: data = 12'h396;
        15'h368E: data = 12'h3A9;
        15'h368F: data = 12'h3C3;
        15'h3690: data = 12'h3D9;
        15'h3691: data = 12'h3ED;
        15'h3692: data = 12'h3FE;
        15'h3693: data = 12'h414;
        15'h3694: data = 12'h42D;
        15'h3695: data = 12'h445;
        15'h3696: data = 12'h455;
        15'h3697: data = 12'h46B;
        15'h3698: data = 12'h483;
        15'h3699: data = 12'h49A;
        15'h369A: data = 12'h4AC;
        15'h369B: data = 12'h4BC;
        15'h369C: data = 12'h4CC;
        15'h369D: data = 12'h4DF;
        15'h369E: data = 12'h4F7;
        15'h369F: data = 12'h50A;
        15'h36A0: data = 12'h517;
        15'h36A1: data = 12'h52C;
        15'h36A2: data = 12'h53D;
        15'h36A3: data = 12'h54D;
        15'h36A4: data = 12'h55E;
        15'h36A5: data = 12'h571;
        15'h36A6: data = 12'h584;
        15'h36A7: data = 12'h594;
        15'h36A8: data = 12'h5A8;
        15'h36A9: data = 12'h5BA;
        15'h36AA: data = 12'h5C7;
        15'h36AB: data = 12'h5D3;
        15'h36AC: data = 12'h5E9;
        15'h36AD: data = 12'h5FC;
        15'h36AE: data = 12'h60A;
        15'h36AF: data = 12'h61B;
        15'h36B0: data = 12'h62B;
        15'h36B1: data = 12'h63D;
        15'h36B2: data = 12'h64F;
        15'h36B3: data = 12'h660;
        15'h36B4: data = 12'h670;
        15'h36B5: data = 12'h67E;
        15'h36B6: data = 12'h68E;
        15'h36B7: data = 12'h6A2;
        15'h36B8: data = 12'h6AF;
        15'h36B9: data = 12'h6C1;
        15'h36BA: data = 12'h6CD;
        15'h36BB: data = 12'h6D4;
        15'h36BC: data = 12'h6E5;
        15'h36BD: data = 12'h6F9;
        15'h36BE: data = 12'h705;
        15'h36BF: data = 12'h70F;
        15'h36C0: data = 12'h721;
        15'h36C1: data = 12'h733;
        15'h36C2: data = 12'h737;
        15'h36C3: data = 12'h745;
        15'h36C4: data = 12'h750;
        15'h36C5: data = 12'h75E;
        15'h36C6: data = 12'h765;
        15'h36C7: data = 12'h777;
        15'h36C8: data = 12'h77C;
        15'h36C9: data = 12'h78F;
        15'h36CA: data = 12'h798;
        15'h36CB: data = 12'h79C;
        15'h36CC: data = 12'h7A5;
        15'h36CD: data = 12'h7B2;
        15'h36CE: data = 12'h7B9;
        15'h36CF: data = 12'h7C3;
        15'h36D0: data = 12'h7C7;
        15'h36D1: data = 12'h7D0;
        15'h36D2: data = 12'h7D5;
        15'h36D3: data = 12'h7E1;
        15'h36D4: data = 12'h7E9;
        15'h36D5: data = 12'h7EF;
        15'h36D6: data = 12'h7F6;
        15'h36D7: data = 12'h7FB;
        15'h36D8: data = 12'h803;
        15'h36D9: data = 12'h808;
        15'h36DA: data = 12'h80C;
        15'h36DB: data = 12'h812;
        15'h36DC: data = 12'h082;
        15'h36DD: data = 12'h092;
        15'h36DE: data = 12'h09B;
        15'h36DF: data = 12'h09C;
        15'h36E0: data = 12'h09E;
        15'h36E1: data = 12'h0A6;
        15'h36E2: data = 12'h0A5;
        15'h36E3: data = 12'h0AE;
        15'h36E4: data = 12'h0B0;
        15'h36E5: data = 12'h0AF;
        15'h36E6: data = 12'h0B6;
        15'h36E7: data = 12'h0B6;
        15'h36E8: data = 12'h0B6;
        15'h36E9: data = 12'h0B7;
        15'h36EA: data = 12'h0C2;
        15'h36EB: data = 12'h0C3;
        15'h36EC: data = 12'h0C8;
        15'h36ED: data = 12'h0C9;
        15'h36EE: data = 12'h0CC;
        15'h36EF: data = 12'h0D0;
        15'h36F0: data = 12'h0D2;
        15'h36F1: data = 12'h0CF;
        15'h36F2: data = 12'h0CD;
        15'h36F3: data = 12'h0CD;
        15'h36F4: data = 12'h0CC;
        15'h36F5: data = 12'h0C7;
        15'h36F6: data = 12'h0C1;
        15'h36F7: data = 12'h0BF;
        15'h36F8: data = 12'h0B2;
        15'h36F9: data = 12'h0AE;
        15'h36FA: data = 12'h0A4;
        15'h36FB: data = 12'h0A9;
        15'h36FC: data = 12'h0A5;
        15'h36FD: data = 12'h0A8;
        15'h36FE: data = 12'h0A8;
        15'h36FF: data = 12'h0A1;
        15'h3700: data = 12'h0A6;
        15'h3701: data = 12'h09F;
        15'h3702: data = 12'h093;
        15'h3703: data = 12'h089;
        15'h3704: data = 12'h078;
        15'h3705: data = 12'h076;
        15'h3706: data = 12'h06F;
        15'h3707: data = 12'h066;
        15'h3708: data = 12'h064;
        15'h3709: data = 12'h060;
        15'h370A: data = 12'h05F;
        15'h370B: data = 12'h057;
        15'h370C: data = 12'h049;
        15'h370D: data = 12'h483;
        15'h370E: data = 12'h7BB;
        15'h370F: data = 12'h7A7;
        15'h3710: data = 12'h79D;
        15'h3711: data = 12'h78E;
        15'h3712: data = 12'h78B;
        15'h3713: data = 12'h78A;
        15'h3714: data = 12'h77A;
        15'h3715: data = 12'h76E;
        15'h3716: data = 12'h761;
        15'h3717: data = 12'h74F;
        15'h3718: data = 12'h73D;
        15'h3719: data = 12'h72E;
        15'h371A: data = 12'h720;
        15'h371B: data = 12'h717;
        15'h371C: data = 12'h70C;
        15'h371D: data = 12'h707;
        15'h371E: data = 12'h6FC;
        15'h371F: data = 12'h6ED;
        15'h3720: data = 12'h6DF;
        15'h3721: data = 12'h6CF;
        15'h3722: data = 12'h6BB;
        15'h3723: data = 12'h6A7;
        15'h3724: data = 12'h696;
        15'h3725: data = 12'h688;
        15'h3726: data = 12'h677;
        15'h3727: data = 12'h66D;
        15'h3728: data = 12'h665;
        15'h3729: data = 12'h654;
        15'h372A: data = 12'h646;
        15'h372B: data = 12'h635;
        15'h372C: data = 12'h62C;
        15'h372D: data = 12'h615;
        15'h372E: data = 12'h5FF;
        15'h372F: data = 12'h5F1;
        15'h3730: data = 12'h5D0;
        15'h3731: data = 12'h5C1;
        15'h3732: data = 12'h5B0;
        15'h3733: data = 12'h59E;
        15'h3734: data = 12'h58A;
        15'h3735: data = 12'h575;
        15'h3736: data = 12'h56D;
        15'h3737: data = 12'h55E;
        15'h3738: data = 12'h54F;
        15'h3739: data = 12'h53F;
        15'h373A: data = 12'h52D;
        15'h373B: data = 12'h517;
        15'h373C: data = 12'h507;
        15'h373D: data = 12'h4F5;
        15'h373E: data = 12'h4DE;
        15'h373F: data = 12'h4C7;
        15'h3740: data = 12'h4B5;
        15'h3741: data = 12'h499;
        15'h3742: data = 12'h485;
        15'h3743: data = 12'h46B;
        15'h3744: data = 12'h455;
        15'h3745: data = 12'h441;
        15'h3746: data = 12'h42B;
        15'h3747: data = 12'h417;
        15'h3748: data = 12'h3FE;
        15'h3749: data = 12'h3E5;
        15'h374A: data = 12'h3D2;
        15'h374B: data = 12'h3BA;
        15'h374C: data = 12'h3AA;
        15'h374D: data = 12'h38B;
        15'h374E: data = 12'h37C;
        15'h374F: data = 12'h369;
        15'h3750: data = 12'h351;
        15'h3751: data = 12'h33B;
        15'h3752: data = 12'h328;
        15'h3753: data = 12'h312;
        15'h3754: data = 12'h2FC;
        15'h3755: data = 12'h2E7;
        15'h3756: data = 12'h2D4;
        15'h3757: data = 12'h2BF;
        15'h3758: data = 12'h2A4;
        15'h3759: data = 12'h28E;
        15'h375A: data = 12'h27F;
        15'h375B: data = 12'h263;
        15'h375C: data = 12'h248;
        15'h375D: data = 12'h232;
        15'h375E: data = 12'h21C;
        15'h375F: data = 12'h208;
        15'h3760: data = 12'h1F3;
        15'h3761: data = 12'h1D9;
        15'h3762: data = 12'h1C2;
        15'h3763: data = 12'h1AB;
        15'h3764: data = 12'h192;
        15'h3765: data = 12'h17E;
        15'h3766: data = 12'h167;
        15'h3767: data = 12'h151;
        15'h3768: data = 12'h139;
        15'h3769: data = 12'h11E;
        15'h376A: data = 12'h109;
        15'h376B: data = 12'h0F5;
        15'h376C: data = 12'h0DA;
        15'h376D: data = 12'h0BE;
        15'h376E: data = 12'h0A6;
        15'h376F: data = 12'h091;
        15'h3770: data = 12'h080;
        15'h3771: data = 12'h066;
        15'h3772: data = 12'h04D;
        15'h3773: data = 12'h7E3;
        15'h3774: data = 12'h7D0;
        15'h3775: data = 12'h7B9;
        15'h3776: data = 12'h7A5;
        15'h3777: data = 12'h78E;
        15'h3778: data = 12'h776;
        15'h3779: data = 12'h75A;
        15'h377A: data = 12'h74E;
        15'h377B: data = 12'h736;
        15'h377C: data = 12'h720;
        15'h377D: data = 12'h706;
        15'h377E: data = 12'h6EC;
        15'h377F: data = 12'h6DD;
        15'h3780: data = 12'h6C7;
        15'h3781: data = 12'h6AE;
        15'h3782: data = 12'h697;
        15'h3783: data = 12'h681;
        15'h3784: data = 12'h668;
        15'h3785: data = 12'h655;
        15'h3786: data = 12'h63C;
        15'h3787: data = 12'h629;
        15'h3788: data = 12'h617;
        15'h3789: data = 12'h5FA;
        15'h378A: data = 12'h5E5;
        15'h378B: data = 12'h5D1;
        15'h378C: data = 12'h5BF;
        15'h378D: data = 12'h5A3;
        15'h378E: data = 12'h58A;
        15'h378F: data = 12'h577;
        15'h3790: data = 12'h564;
        15'h3791: data = 12'h54D;
        15'h3792: data = 12'h537;
        15'h3793: data = 12'h520;
        15'h3794: data = 12'h508;
        15'h3795: data = 12'h4F6;
        15'h3796: data = 12'h4E1;
        15'h3797: data = 12'h4CA;
        15'h3798: data = 12'h4B5;
        15'h3799: data = 12'h4A3;
        15'h379A: data = 12'h48F;
        15'h379B: data = 12'h47C;
        15'h379C: data = 12'h467;
        15'h379D: data = 12'h455;
        15'h379E: data = 12'h445;
        15'h379F: data = 12'h432;
        15'h37A0: data = 12'h424;
        15'h37A1: data = 12'h412;
        15'h37A2: data = 12'h402;
        15'h37A3: data = 12'h3F5;
        15'h37A4: data = 12'h3E7;
        15'h37A5: data = 12'h3D0;
        15'h37A6: data = 12'h3C4;
        15'h37A7: data = 12'h3B1;
        15'h37A8: data = 12'h39D;
        15'h37A9: data = 12'h395;
        15'h37AA: data = 12'h379;
        15'h37AB: data = 12'h368;
        15'h37AC: data = 12'h359;
        15'h37AD: data = 12'h345;
        15'h37AE: data = 12'h335;
        15'h37AF: data = 12'h322;
        15'h37B0: data = 12'h311;
        15'h37B1: data = 12'h2FE;
        15'h37B2: data = 12'h2EE;
        15'h37B3: data = 12'h2DD;
        15'h37B4: data = 12'h2D0;
        15'h37B5: data = 12'h2C8;
        15'h37B6: data = 12'h2BE;
        15'h37B7: data = 12'h2B3;
        15'h37B8: data = 12'h2A7;
        15'h37B9: data = 12'h29C;
        15'h37BA: data = 12'h295;
        15'h37BB: data = 12'h287;
        15'h37BC: data = 12'h280;
        15'h37BD: data = 12'h26D;
        15'h37BE: data = 12'h264;
        15'h37BF: data = 12'h253;
        15'h37C0: data = 12'h249;
        15'h37C1: data = 12'h235;
        15'h37C2: data = 12'h226;
        15'h37C3: data = 12'h217;
        15'h37C4: data = 12'h20C;
        15'h37C5: data = 12'h206;
        15'h37C6: data = 12'h200;
        15'h37C7: data = 12'h1F2;
        15'h37C8: data = 12'h1F0;
        15'h37C9: data = 12'h1EC;
        15'h37CA: data = 12'h1EA;
        15'h37CB: data = 12'h1DE;
        15'h37CC: data = 12'h1D7;
        15'h37CD: data = 12'h1CA;
        15'h37CE: data = 12'h1C2;
        15'h37CF: data = 12'h1C3;
        15'h37D0: data = 12'h1B6;
        15'h37D1: data = 12'h1A6;
        15'h37D2: data = 12'h19D;
        15'h37D3: data = 12'h194;
        15'h37D4: data = 12'h18F;
        15'h37D5: data = 12'h18C;
        15'h37D6: data = 12'h184;
        15'h37D7: data = 12'h181;
        15'h37D8: data = 12'h185;
        15'h37D9: data = 12'h183;
        15'h37DA: data = 12'h184;
        15'h37DB: data = 12'h17E;
        15'h37DC: data = 12'h17F;
        15'h37DD: data = 12'h174;
        15'h37DE: data = 12'h173;
        15'h37DF: data = 12'h173;
        15'h37E0: data = 12'h168;
        15'h37E1: data = 12'h163;
        15'h37E2: data = 12'h162;
        15'h37E3: data = 12'h15F;
        15'h37E4: data = 12'h154;
        15'h37E5: data = 12'h157;
        15'h37E6: data = 12'h157;
        15'h37E7: data = 12'h15B;
        15'h37E8: data = 12'h15E;
        15'h37E9: data = 12'h166;
        15'h37EA: data = 12'h166;
        15'h37EB: data = 12'h16F;
        15'h37EC: data = 12'h173;
        15'h37ED: data = 12'h16F;
        15'h37EE: data = 12'h16D;
        15'h37EF: data = 12'h16C;
        15'h37F0: data = 12'h171;
        15'h37F1: data = 12'h16D;
        15'h37F2: data = 12'h16E;
        15'h37F3: data = 12'h16B;
        15'h37F4: data = 12'h170;
        15'h37F5: data = 12'h174;
        15'h37F6: data = 12'h17A;
        15'h37F7: data = 12'h17F;
        15'h37F8: data = 12'h18B;
        15'h37F9: data = 12'h18F;
        15'h37FA: data = 12'h19A;
        15'h37FB: data = 12'h1A3;
        15'h37FC: data = 12'h1AE;
        15'h37FD: data = 12'h1B6;
        15'h37FE: data = 12'h1B6;
        15'h37FF: data = 12'h1BA;
        15'h3800: data = 12'h1BE;
        15'h3801: data = 12'h1C4;
        15'h3802: data = 12'h1CA;
        15'h3803: data = 12'h1CB;
        15'h3804: data = 12'h1D1;
        15'h3805: data = 12'h1D9;
        15'h3806: data = 12'h1E0;
        15'h3807: data = 12'h1EF;
        15'h3808: data = 12'h1F9;
        15'h3809: data = 12'h202;
        15'h380A: data = 12'h215;
        15'h380B: data = 12'h21C;
        15'h380C: data = 12'h232;
        15'h380D: data = 12'h238;
        15'h380E: data = 12'h24A;
        15'h380F: data = 12'h24E;
        15'h3810: data = 12'h25D;
        15'h3811: data = 12'h264;
        15'h3812: data = 12'h273;
        15'h3813: data = 12'h27A;
        15'h3814: data = 12'h283;
        15'h3815: data = 12'h28E;
        15'h3816: data = 12'h293;
        15'h3817: data = 12'h2A3;
        15'h3818: data = 12'h2B0;
        15'h3819: data = 12'h2C0;
        15'h381A: data = 12'h2CF;
        15'h381B: data = 12'h2DC;
        15'h381C: data = 12'h2EF;
        15'h381D: data = 12'h301;
        15'h381E: data = 12'h310;
        15'h381F: data = 12'h322;
        15'h3820: data = 12'h337;
        15'h3821: data = 12'h347;
        15'h3822: data = 12'h358;
        15'h3823: data = 12'h364;
        15'h3824: data = 12'h375;
        15'h3825: data = 12'h382;
        15'h3826: data = 12'h397;
        15'h3827: data = 12'h39D;
        15'h3828: data = 12'h3B1;
        15'h3829: data = 12'h3BA;
        15'h382A: data = 12'h3CB;
        15'h382B: data = 12'h3DD;
        15'h382C: data = 12'h3ED;
        15'h382D: data = 12'h3FA;
        15'h382E: data = 12'h413;
        15'h382F: data = 12'h423;
        15'h3830: data = 12'h43B;
        15'h3831: data = 12'h451;
        15'h3832: data = 12'h466;
        15'h3833: data = 12'h47B;
        15'h3834: data = 12'h490;
        15'h3835: data = 12'h4A7;
        15'h3836: data = 12'h4B8;
        15'h3837: data = 12'h4D0;
        15'h3838: data = 12'h4E6;
        15'h3839: data = 12'h4FB;
        15'h383A: data = 12'h50C;
        15'h383B: data = 12'h520;
        15'h383C: data = 12'h52E;
        15'h383D: data = 12'h545;
        15'h383E: data = 12'h55A;
        15'h383F: data = 12'h569;
        15'h3840: data = 12'h579;
        15'h3841: data = 12'h58A;
        15'h3842: data = 12'h5A4;
        15'h3843: data = 12'h5B9;
        15'h3844: data = 12'h5CB;
        15'h3845: data = 12'h5E4;
        15'h3846: data = 12'h5FB;
        15'h3847: data = 12'h615;
        15'h3848: data = 12'h62D;
        15'h3849: data = 12'h645;
        15'h384A: data = 12'h661;
        15'h384B: data = 12'h674;
        15'h384C: data = 12'h691;
        15'h384D: data = 12'h6A2;
        15'h384E: data = 12'h6BA;
        15'h384F: data = 12'h6D2;
        15'h3850: data = 12'h6E4;
        15'h3851: data = 12'h6FC;
        15'h3852: data = 12'h711;
        15'h3853: data = 12'h722;
        15'h3854: data = 12'h73A;
        15'h3855: data = 12'h74A;
        15'h3856: data = 12'h75F;
        15'h3857: data = 12'h776;
        15'h3858: data = 12'h790;
        15'h3859: data = 12'h7A0;
        15'h385A: data = 12'h7B9;
        15'h385B: data = 12'h7D3;
        15'h385C: data = 12'h7E8;
        15'h385D: data = 12'h800;
        15'h385E: data = 12'h06F;
        15'h385F: data = 12'h088;
        15'h3860: data = 12'h09F;
        15'h3861: data = 12'h0B5;
        15'h3862: data = 12'h0D0;
        15'h3863: data = 12'h0E9;
        15'h3864: data = 12'h102;
        15'h3865: data = 12'h117;
        15'h3866: data = 12'h12D;
        15'h3867: data = 12'h147;
        15'h3868: data = 12'h158;
        15'h3869: data = 12'h16E;
        15'h386A: data = 12'h187;
        15'h386B: data = 12'h19D;
        15'h386C: data = 12'h1B5;
        15'h386D: data = 12'h1C4;
        15'h386E: data = 12'h1DC;
        15'h386F: data = 12'h1F2;
        15'h3870: data = 12'h207;
        15'h3871: data = 12'h21C;
        15'h3872: data = 12'h234;
        15'h3873: data = 12'h24C;
        15'h3874: data = 12'h262;
        15'h3875: data = 12'h276;
        15'h3876: data = 12'h289;
        15'h3877: data = 12'h2A2;
        15'h3878: data = 12'h2BC;
        15'h3879: data = 12'h2D1;
        15'h387A: data = 12'h2EB;
        15'h387B: data = 12'h306;
        15'h387C: data = 12'h321;
        15'h387D: data = 12'h32F;
        15'h387E: data = 12'h348;
        15'h387F: data = 12'h366;
        15'h3880: data = 12'h379;
        15'h3881: data = 12'h39A;
        15'h3882: data = 12'h3A9;
        15'h3883: data = 12'h3C1;
        15'h3884: data = 12'h3DD;
        15'h3885: data = 12'h3F0;
        15'h3886: data = 12'h400;
        15'h3887: data = 12'h41A;
        15'h3888: data = 12'h42F;
        15'h3889: data = 12'h446;
        15'h388A: data = 12'h456;
        15'h388B: data = 12'h469;
        15'h388C: data = 12'h482;
        15'h388D: data = 12'h498;
        15'h388E: data = 12'h4AC;
        15'h388F: data = 12'h4BB;
        15'h3890: data = 12'h4CB;
        15'h3891: data = 12'h4DD;
        15'h3892: data = 12'h4F6;
        15'h3893: data = 12'h508;
        15'h3894: data = 12'h519;
        15'h3895: data = 12'h52C;
        15'h3896: data = 12'h53D;
        15'h3897: data = 12'h54A;
        15'h3898: data = 12'h55D;
        15'h3899: data = 12'h56B;
        15'h389A: data = 12'h583;
        15'h389B: data = 12'h594;
        15'h389C: data = 12'h5A5;
        15'h389D: data = 12'h5B7;
        15'h389E: data = 12'h5C8;
        15'h389F: data = 12'h5D3;
        15'h38A0: data = 12'h5E9;
        15'h38A1: data = 12'h5F8;
        15'h38A2: data = 12'h60B;
        15'h38A3: data = 12'h61A;
        15'h38A4: data = 12'h62A;
        15'h38A5: data = 12'h63B;
        15'h38A6: data = 12'h650;
        15'h38A7: data = 12'h65E;
        15'h38A8: data = 12'h66D;
        15'h38A9: data = 12'h67E;
        15'h38AA: data = 12'h68F;
        15'h38AB: data = 12'h6A0;
        15'h38AC: data = 12'h6AE;
        15'h38AD: data = 12'h6BD;
        15'h38AE: data = 12'h6D0;
        15'h38AF: data = 12'h6D7;
        15'h38B0: data = 12'h6E9;
        15'h38B1: data = 12'h6F9;
        15'h38B2: data = 12'h707;
        15'h38B3: data = 12'h712;
        15'h38B4: data = 12'h721;
        15'h38B5: data = 12'h731;
        15'h38B6: data = 12'h739;
        15'h38B7: data = 12'h745;
        15'h38B8: data = 12'h74C;
        15'h38B9: data = 12'h75F;
        15'h38BA: data = 12'h765;
        15'h38BB: data = 12'h777;
        15'h38BC: data = 12'h77C;
        15'h38BD: data = 12'h78D;
        15'h38BE: data = 12'h795;
        15'h38BF: data = 12'h79D;
        15'h38C0: data = 12'h7A6;
        15'h38C1: data = 12'h7B0;
        15'h38C2: data = 12'h7BB;
        15'h38C3: data = 12'h7BD;
        15'h38C4: data = 12'h7C6;
        15'h38C5: data = 12'h7CE;
        15'h38C6: data = 12'h7D7;
        15'h38C7: data = 12'h7E0;
        15'h38C8: data = 12'h7EB;
        15'h38C9: data = 12'h7F0;
        15'h38CA: data = 12'h7F7;
        15'h38CB: data = 12'h7FD;
        15'h38CC: data = 12'h801;
        15'h38CD: data = 12'h807;
        15'h38CE: data = 12'h805;
        15'h38CF: data = 12'h80F;
        15'h38D0: data = 12'h887;
        15'h38D1: data = 12'h08B;
        15'h38D2: data = 12'h097;
        15'h38D3: data = 12'h096;
        15'h38D4: data = 12'h09B;
        15'h38D5: data = 12'h0A0;
        15'h38D6: data = 12'h0A7;
        15'h38D7: data = 12'h0AA;
        15'h38D8: data = 12'h0AF;
        15'h38D9: data = 12'h0AB;
        15'h38DA: data = 12'h0B6;
        15'h38DB: data = 12'h0B7;
        15'h38DC: data = 12'h0B6;
        15'h38DD: data = 12'h0B7;
        15'h38DE: data = 12'h0C2;
        15'h38DF: data = 12'h0C4;
        15'h38E0: data = 12'h0CA;
        15'h38E1: data = 12'h0CC;
        15'h38E2: data = 12'h0CE;
        15'h38E3: data = 12'h0D0;
        15'h38E4: data = 12'h0D3;
        15'h38E5: data = 12'h0CB;
        15'h38E6: data = 12'h0CC;
        15'h38E7: data = 12'h0CA;
        15'h38E8: data = 12'h0CA;
        15'h38E9: data = 12'h0C6;
        15'h38EA: data = 12'h0BB;
        15'h38EB: data = 12'h0BA;
        15'h38EC: data = 12'h0A9;
        15'h38ED: data = 12'h0AC;
        15'h38EE: data = 12'h0A1;
        15'h38EF: data = 12'h0A7;
        15'h38F0: data = 12'h0A4;
        15'h38F1: data = 12'h0AD;
        15'h38F2: data = 12'h0A9;
        15'h38F3: data = 12'h0A5;
        15'h38F4: data = 12'h0A8;
        15'h38F5: data = 12'h09D;
        15'h38F6: data = 12'h093;
        15'h38F7: data = 12'h084;
        15'h38F8: data = 12'h074;
        15'h38F9: data = 12'h076;
        15'h38FA: data = 12'h06D;
        15'h38FB: data = 12'h067;
        15'h38FC: data = 12'h064;
        15'h38FD: data = 12'h065;
        15'h38FE: data = 12'h060;
        15'h38FF: data = 12'h054;
        15'h3900: data = 12'h049;
        15'h3901: data = 12'h7C7;
        15'h3902: data = 12'h7B6;
        15'h3903: data = 12'h7A6;
        15'h3904: data = 12'h79F;
        15'h3905: data = 12'h791;
        15'h3906: data = 12'h78C;
        15'h3907: data = 12'h786;
        15'h3908: data = 12'h77C;
        15'h3909: data = 12'h76D;
        15'h390A: data = 12'h75D;
        15'h390B: data = 12'h74D;
        15'h390C: data = 12'h73A;
        15'h390D: data = 12'h72E;
        15'h390E: data = 12'h724;
        15'h390F: data = 12'h716;
        15'h3910: data = 12'h70C;
        15'h3911: data = 12'h706;
        15'h3912: data = 12'h6FA;
        15'h3913: data = 12'h6EE;
        15'h3914: data = 12'h6DE;
        15'h3915: data = 12'h6CE;
        15'h3916: data = 12'h6B9;
        15'h3917: data = 12'h6A8;
        15'h3918: data = 12'h695;
        15'h3919: data = 12'h686;
        15'h391A: data = 12'h678;
        15'h391B: data = 12'h66D;
        15'h391C: data = 12'h661;
        15'h391D: data = 12'h653;
        15'h391E: data = 12'h643;
        15'h391F: data = 12'h635;
        15'h3920: data = 12'h629;
        15'h3921: data = 12'h613;
        15'h3922: data = 12'h601;
        15'h3923: data = 12'h5EE;
        15'h3924: data = 12'h5D0;
        15'h3925: data = 12'h5BF;
        15'h3926: data = 12'h5AF;
        15'h3927: data = 12'h59B;
        15'h3928: data = 12'h588;
        15'h3929: data = 12'h578;
        15'h392A: data = 12'h56B;
        15'h392B: data = 12'h55D;
        15'h392C: data = 12'h551;
        15'h392D: data = 12'h53F;
        15'h392E: data = 12'h52A;
        15'h392F: data = 12'h519;
        15'h3930: data = 12'h506;
        15'h3931: data = 12'h4F7;
        15'h3932: data = 12'h4DC;
        15'h3933: data = 12'h4C7;
        15'h3934: data = 12'h4B7;
        15'h3935: data = 12'h49B;
        15'h3936: data = 12'h485;
        15'h3937: data = 12'h46C;
        15'h3938: data = 12'h458;
        15'h3939: data = 12'h441;
        15'h393A: data = 12'h42A;
        15'h393B: data = 12'h415;
        15'h393C: data = 12'h3FF;
        15'h393D: data = 12'h3E2;
        15'h393E: data = 12'h3CE;
        15'h393F: data = 12'h3BC;
        15'h3940: data = 12'h3A8;
        15'h3941: data = 12'h38E;
        15'h3942: data = 12'h37A;
        15'h3943: data = 12'h367;
        15'h3944: data = 12'h34E;
        15'h3945: data = 12'h33A;
        15'h3946: data = 12'h323;
        15'h3947: data = 12'h30F;
        15'h3948: data = 12'h2F7;
        15'h3949: data = 12'h2E2;
        15'h394A: data = 12'h2CF;
        15'h394B: data = 12'h2BE;
        15'h394C: data = 12'h2A3;
        15'h394D: data = 12'h286;
        15'h394E: data = 12'h27B;
        15'h394F: data = 12'h260;
        15'h3950: data = 12'h245;
        15'h3951: data = 12'h232;
        15'h3952: data = 12'h217;
        15'h3953: data = 12'h205;
        15'h3954: data = 12'h1EC;
        15'h3955: data = 12'h1D5;
        15'h3956: data = 12'h1BE;
        15'h3957: data = 12'h1AA;
        15'h3958: data = 12'h191;
        15'h3959: data = 12'h17C;
        15'h395A: data = 12'h165;
        15'h395B: data = 12'h14F;
        15'h395C: data = 12'h137;
        15'h395D: data = 12'h11A;
        15'h395E: data = 12'h107;
        15'h395F: data = 12'h0F2;
        15'h3960: data = 12'h0D8;
        15'h3961: data = 12'h0BF;
        15'h3962: data = 12'h0A6;
        15'h3963: data = 12'h090;
        15'h3964: data = 12'h07C;
        15'h3965: data = 12'h064;
        15'h3966: data = 12'h04B;
        15'h3967: data = 12'h7E2;
        15'h3968: data = 12'h7CD;
        15'h3969: data = 12'h7B6;
        15'h396A: data = 12'h7A3;
        15'h396B: data = 12'h78E;
        15'h396C: data = 12'h774;
        15'h396D: data = 12'h758;
        15'h396E: data = 12'h749;
        15'h396F: data = 12'h735;
        15'h3970: data = 12'h71C;
        15'h3971: data = 12'h706;
        15'h3972: data = 12'h6EB;
        15'h3973: data = 12'h6DA;
        15'h3974: data = 12'h6C5;
        15'h3975: data = 12'h6B0;
        15'h3976: data = 12'h694;
        15'h3977: data = 12'h683;
        15'h3978: data = 12'h66A;
        15'h3979: data = 12'h655;
        15'h397A: data = 12'h63C;
        15'h397B: data = 12'h62A;
        15'h397C: data = 12'h615;
        15'h397D: data = 12'h5F9;
        15'h397E: data = 12'h5E5;
        15'h397F: data = 12'h5D1;
        15'h3980: data = 12'h5BC;
        15'h3981: data = 12'h5A1;
        15'h3982: data = 12'h58A;
        15'h3983: data = 12'h577;
        15'h3984: data = 12'h562;
        15'h3985: data = 12'h54D;
        15'h3986: data = 12'h539;
        15'h3987: data = 12'h522;
        15'h3988: data = 12'h50E;
        15'h3989: data = 12'h4F8;
        15'h398A: data = 12'h4DE;
        15'h398B: data = 12'h4CB;
        15'h398C: data = 12'h4B4;
        15'h398D: data = 12'h4A3;
        15'h398E: data = 12'h48F;
        15'h398F: data = 12'h476;
        15'h3990: data = 12'h464;
        15'h3991: data = 12'h454;
        15'h3992: data = 12'h442;
        15'h3993: data = 12'h432;
        15'h3994: data = 12'h422;
        15'h3995: data = 12'h40C;
        15'h3996: data = 12'h401;
        15'h3997: data = 12'h3F4;
        15'h3998: data = 12'h3E6;
        15'h3999: data = 12'h3D1;
        15'h399A: data = 12'h3C1;
        15'h399B: data = 12'h3AE;
        15'h399C: data = 12'h39D;
        15'h399D: data = 12'h393;
        15'h399E: data = 12'h378;
        15'h399F: data = 12'h367;
        15'h39A0: data = 12'h355;
        15'h39A1: data = 12'h344;
        15'h39A2: data = 12'h333;
        15'h39A3: data = 12'h31F;
        15'h39A4: data = 12'h310;
        15'h39A5: data = 12'h2FE;
        15'h39A6: data = 12'h2EE;
        15'h39A7: data = 12'h2DD;
        15'h39A8: data = 12'h2CD;
        15'h39A9: data = 12'h2CD;
        15'h39AA: data = 12'h2BF;
        15'h39AB: data = 12'h2B5;
        15'h39AC: data = 12'h2AA;
        15'h39AD: data = 12'h29B;
        15'h39AE: data = 12'h293;
        15'h39AF: data = 12'h285;
        15'h39B0: data = 12'h27A;
        15'h39B1: data = 12'h26C;
        15'h39B2: data = 12'h264;
        15'h39B3: data = 12'h252;
        15'h39B4: data = 12'h246;
        15'h39B5: data = 12'h230;
        15'h39B6: data = 12'h223;
        15'h39B7: data = 12'h213;
        15'h39B8: data = 12'h20C;
        15'h39B9: data = 12'h209;
        15'h39BA: data = 12'h203;
        15'h39BB: data = 12'h1F6;
        15'h39BC: data = 12'h1F2;
        15'h39BD: data = 12'h1EC;
        15'h39BE: data = 12'h1E9;
        15'h39BF: data = 12'h1E4;
        15'h39C0: data = 12'h1D4;
        15'h39C1: data = 12'h1C9;
        15'h39C2: data = 12'h1C0;
        15'h39C3: data = 12'h1C0;
        15'h39C4: data = 12'h1B8;
        15'h39C5: data = 12'h1A6;
        15'h39C6: data = 12'h19D;
        15'h39C7: data = 12'h193;
        15'h39C8: data = 12'h191;
        15'h39C9: data = 12'h18A;
        15'h39CA: data = 12'h185;
        15'h39CB: data = 12'h185;
        15'h39CC: data = 12'h185;
        15'h39CD: data = 12'h184;
        15'h39CE: data = 12'h186;
        15'h39CF: data = 12'h180;
        15'h39D0: data = 12'h17F;
        15'h39D1: data = 12'h177;
        15'h39D2: data = 12'h175;
        15'h39D3: data = 12'h174;
        15'h39D4: data = 12'h166;
        15'h39D5: data = 12'h161;
        15'h39D6: data = 12'h15D;
        15'h39D7: data = 12'h15E;
        15'h39D8: data = 12'h156;
        15'h39D9: data = 12'h155;
        15'h39DA: data = 12'h159;
        15'h39DB: data = 12'h15C;
        15'h39DC: data = 12'h164;
        15'h39DD: data = 12'h163;
        15'h39DE: data = 12'h167;
        15'h39DF: data = 12'h16F;
        15'h39E0: data = 12'h16F;
        15'h39E1: data = 12'h16D;
        15'h39E2: data = 12'h16E;
        15'h39E3: data = 12'h16C;
        15'h39E4: data = 12'h171;
        15'h39E5: data = 12'h16B;
        15'h39E6: data = 12'h16D;
        15'h39E7: data = 12'h16C;
        15'h39E8: data = 12'h16D;
        15'h39E9: data = 12'h174;
        15'h39EA: data = 12'h17C;
        15'h39EB: data = 12'h183;
        15'h39EC: data = 12'h18C;
        15'h39ED: data = 12'h18F;
        15'h39EE: data = 12'h19D;
        15'h39EF: data = 12'h1A3;
        15'h39F0: data = 12'h1AE;
        15'h39F1: data = 12'h1B1;
        15'h39F2: data = 12'h1B4;
        15'h39F3: data = 12'h1B8;
        15'h39F4: data = 12'h1C0;
        15'h39F5: data = 12'h1C3;
        15'h39F6: data = 12'h1C7;
        15'h39F7: data = 12'h1C8;
        15'h39F8: data = 12'h1D1;
        15'h39F9: data = 12'h1D7;
        15'h39FA: data = 12'h1E0;
        15'h39FB: data = 12'h1ED;
        15'h39FC: data = 12'h1F7;
        15'h39FD: data = 12'h206;
        15'h39FE: data = 12'h219;
        15'h39FF: data = 12'h21C;
        15'h3A00: data = 12'h22E;
        15'h3A01: data = 12'h238;
        15'h3A02: data = 12'h247;
        15'h3A03: data = 12'h24D;
        15'h3A04: data = 12'h25D;
        15'h3A05: data = 12'h26A;
        15'h3A06: data = 12'h272;
        15'h3A07: data = 12'h278;
        15'h3A08: data = 12'h284;
        15'h3A09: data = 12'h28B;
        15'h3A0A: data = 12'h292;
        15'h3A0B: data = 12'h2A2;
        15'h3A0C: data = 12'h2AF;
        15'h3A0D: data = 12'h2BD;
        15'h3A0E: data = 12'h2CF;
        15'h3A0F: data = 12'h2D9;
        15'h3A10: data = 12'h2ED;
        15'h3A11: data = 12'h2FF;
        15'h3A12: data = 12'h314;
        15'h3A13: data = 12'h325;
        15'h3A14: data = 12'h336;
        15'h3A15: data = 12'h346;
        15'h3A16: data = 12'h356;
        15'h3A17: data = 12'h368;
        15'h3A18: data = 12'h375;
        15'h3A19: data = 12'h383;
        15'h3A1A: data = 12'h397;
        15'h3A1B: data = 12'h39D;
        15'h3A1C: data = 12'h3B1;
        15'h3A1D: data = 12'h3BB;
        15'h3A1E: data = 12'h3C9;
        15'h3A1F: data = 12'h3DF;
        15'h3A20: data = 12'h3ED;
        15'h3A21: data = 12'h3FC;
        15'h3A22: data = 12'h418;
        15'h3A23: data = 12'h425;
        15'h3A24: data = 12'h43B;
        15'h3A25: data = 12'h451;
        15'h3A26: data = 12'h462;
        15'h3A27: data = 12'h47E;
        15'h3A28: data = 12'h493;
        15'h3A29: data = 12'h4AA;
        15'h3A2A: data = 12'h4B8;
        15'h3A2B: data = 12'h4CF;
        15'h3A2C: data = 12'h4E6;
        15'h3A2D: data = 12'h4F9;
        15'h3A2E: data = 12'h50D;
        15'h3A2F: data = 12'h51E;
        15'h3A30: data = 12'h52F;
        15'h3A31: data = 12'h546;
        15'h3A32: data = 12'h557;
        15'h3A33: data = 12'h569;
        15'h3A34: data = 12'h57A;
        15'h3A35: data = 12'h58C;
        15'h3A36: data = 12'h5A2;
        15'h3A37: data = 12'h5B6;
        15'h3A38: data = 12'h5C8;
        15'h3A39: data = 12'h5E3;
        15'h3A3A: data = 12'h5FA;
        15'h3A3B: data = 12'h611;
        15'h3A3C: data = 12'h62B;
        15'h3A3D: data = 12'h643;
        15'h3A3E: data = 12'h660;
        15'h3A3F: data = 12'h679;
        15'h3A40: data = 12'h690;
        15'h3A41: data = 12'h6A2;
        15'h3A42: data = 12'h6BB;
        15'h3A43: data = 12'h6D3;
        15'h3A44: data = 12'h6E6;
        15'h3A45: data = 12'h6F9;
        15'h3A46: data = 12'h70F;
        15'h3A47: data = 12'h726;
        15'h3A48: data = 12'h741;
        15'h3A49: data = 12'h74D;
        15'h3A4A: data = 12'h761;
        15'h3A4B: data = 12'h776;
        15'h3A4C: data = 12'h791;
        15'h3A4D: data = 12'h7A2;
        15'h3A4E: data = 12'h7B8;
        15'h3A4F: data = 12'h7D4;
        15'h3A50: data = 12'h7E6;
        15'h3A51: data = 12'h7FE;
        15'h3A52: data = 12'h06E;
        15'h3A53: data = 12'h084;
        15'h3A54: data = 12'h099;
        15'h3A55: data = 12'h0B2;
        15'h3A56: data = 12'h0CE;
        15'h3A57: data = 12'h0E7;
        15'h3A58: data = 12'h102;
        15'h3A59: data = 12'h114;
        15'h3A5A: data = 12'h12E;
        15'h3A5B: data = 12'h147;
        15'h3A5C: data = 12'h158;
        15'h3A5D: data = 12'h16F;
        15'h3A5E: data = 12'h183;
        15'h3A5F: data = 12'h19D;
        15'h3A60: data = 12'h1B7;
        15'h3A61: data = 12'h1C5;
        15'h3A62: data = 12'h1DF;
        15'h3A63: data = 12'h1F3;
        15'h3A64: data = 12'h208;
        15'h3A65: data = 12'h21D;
        15'h3A66: data = 12'h234;
        15'h3A67: data = 12'h24C;
        15'h3A68: data = 12'h260;
        15'h3A69: data = 12'h277;
        15'h3A6A: data = 12'h288;
        15'h3A6B: data = 12'h2A6;
        15'h3A6C: data = 12'h2BA;
        15'h3A6D: data = 12'h2D1;
        15'h3A6E: data = 12'h2EA;
        15'h3A6F: data = 12'h303;
        15'h3A70: data = 12'h31E;
        15'h3A71: data = 12'h332;
        15'h3A72: data = 12'h348;
        15'h3A73: data = 12'h365;
        15'h3A74: data = 12'h37B;
        15'h3A75: data = 12'h395;
        15'h3A76: data = 12'h3A9;
        15'h3A77: data = 12'h3C3;
        15'h3A78: data = 12'h3D7;
        15'h3A79: data = 12'h3F1;
        15'h3A7A: data = 12'h401;
        15'h3A7B: data = 12'h416;
        15'h3A7C: data = 12'h42D;
        15'h3A7D: data = 12'h446;
        15'h3A7E: data = 12'h454;
        15'h3A7F: data = 12'h46A;
        15'h3A80: data = 12'h480;
        15'h3A81: data = 12'h498;
        15'h3A82: data = 12'h4AC;
        15'h3A83: data = 12'h4BE;
        15'h3A84: data = 12'h4CF;
        15'h3A85: data = 12'h4E0;
        15'h3A86: data = 12'h4F7;
        15'h3A87: data = 12'h50B;
        15'h3A88: data = 12'h517;
        15'h3A89: data = 12'h52D;
        15'h3A8A: data = 12'h53C;
        15'h3A8B: data = 12'h54C;
        15'h3A8C: data = 12'h560;
        15'h3A8D: data = 12'h570;
        15'h3A8E: data = 12'h587;
        15'h3A8F: data = 12'h594;
        15'h3A90: data = 12'h5A6;
        15'h3A91: data = 12'h5B7;
        15'h3A92: data = 12'h5C7;
        15'h3A93: data = 12'h5D3;
        15'h3A94: data = 12'h5EC;
        15'h3A95: data = 12'h5FB;
        15'h3A96: data = 12'h609;
        15'h3A97: data = 12'h61A;
        15'h3A98: data = 12'h629;
        15'h3A99: data = 12'h638;
        15'h3A9A: data = 12'h64C;
        15'h3A9B: data = 12'h65F;
        15'h3A9C: data = 12'h66D;
        15'h3A9D: data = 12'h67B;
        15'h3A9E: data = 12'h68E;
        15'h3A9F: data = 12'h69D;
        15'h3AA0: data = 12'h6AE;
        15'h3AA1: data = 12'h6BD;
        15'h3AA2: data = 12'h6CB;
        15'h3AA3: data = 12'h6D5;
        15'h3AA4: data = 12'h6E6;
        15'h3AA5: data = 12'h6F6;
        15'h3AA6: data = 12'h705;
        15'h3AA7: data = 12'h713;
        15'h3AA8: data = 12'h721;
        15'h3AA9: data = 12'h731;
        15'h3AAA: data = 12'h738;
        15'h3AAB: data = 12'h743;
        15'h3AAC: data = 12'h74B;
        15'h3AAD: data = 12'h75A;
        15'h3AAE: data = 12'h768;
        15'h3AAF: data = 12'h777;
        15'h3AB0: data = 12'h77D;
        15'h3AB1: data = 12'h790;
        15'h3AB2: data = 12'h794;
        15'h3AB3: data = 12'h79D;
        15'h3AB4: data = 12'h7A5;
        15'h3AB5: data = 12'h7B4;
        15'h3AB6: data = 12'h7BB;
        15'h3AB7: data = 12'h7C1;
        15'h3AB8: data = 12'h7C8;
        15'h3AB9: data = 12'h7D0;
        15'h3ABA: data = 12'h7D6;
        15'h3ABB: data = 12'h7E4;
        15'h3ABC: data = 12'h7EB;
        15'h3ABD: data = 12'h7F1;
        15'h3ABE: data = 12'h7F5;
        15'h3ABF: data = 12'h7FE;
        15'h3AC0: data = 12'h805;
        15'h3AC1: data = 12'h808;
        15'h3AC2: data = 12'h809;
        15'h3AC3: data = 12'h07A;
        15'h3AC4: data = 12'h094;
        15'h3AC5: data = 12'h093;
        15'h3AC6: data = 12'h09D;
        15'h3AC7: data = 12'h0A0;
        15'h3AC8: data = 12'h0A0;
        15'h3AC9: data = 12'h0A6;
        15'h3ACA: data = 12'h0A5;
        15'h3ACB: data = 12'h0AC;
        15'h3ACC: data = 12'h0AE;
        15'h3ACD: data = 12'h0AD;
        15'h3ACE: data = 12'h0B8;
        15'h3ACF: data = 12'h0B7;
        15'h3AD0: data = 12'h0BB;
        15'h3AD1: data = 12'h0B9;
        15'h3AD2: data = 12'h0C2;
        15'h3AD3: data = 12'h0C5;
        15'h3AD4: data = 12'h0C9;
        15'h3AD5: data = 12'h0C9;
        15'h3AD6: data = 12'h0D2;
        15'h3AD7: data = 12'h0D7;
        15'h3AD8: data = 12'h0D4;
        15'h3AD9: data = 12'h0CD;
        15'h3ADA: data = 12'h0D1;
        15'h3ADB: data = 12'h0CF;
        15'h3ADC: data = 12'h0CD;
        15'h3ADD: data = 12'h0C7;
        15'h3ADE: data = 12'h0BD;
        15'h3ADF: data = 12'h0B9;
        15'h3AE0: data = 12'h0AC;
        15'h3AE1: data = 12'h0AE;
        15'h3AE2: data = 12'h0A4;
        15'h3AE3: data = 12'h0A7;
        15'h3AE4: data = 12'h0A9;
        15'h3AE5: data = 12'h0AE;
        15'h3AE6: data = 12'h0AD;
        15'h3AE7: data = 12'h0A4;
        15'h3AE8: data = 12'h0A8;
        15'h3AE9: data = 12'h09C;
        15'h3AEA: data = 12'h090;
        15'h3AEB: data = 12'h084;
        15'h3AEC: data = 12'h072;
        15'h3AED: data = 12'h074;
        15'h3AEE: data = 12'h06C;
        15'h3AEF: data = 12'h069;
        15'h3AF0: data = 12'h06B;
        15'h3AF1: data = 12'h067;
        15'h3AF2: data = 12'h062;
        15'h3AF3: data = 12'h055;
        15'h3AF4: data = 12'h048;
        15'h3AF5: data = 12'h036;
        15'h3AF6: data = 12'h7B4;
        15'h3AF7: data = 12'h7A9;
        15'h3AF8: data = 12'h7A1;
        15'h3AF9: data = 12'h798;
        15'h3AFA: data = 12'h791;
        15'h3AFB: data = 12'h78C;
        15'h3AFC: data = 12'h780;
        15'h3AFD: data = 12'h76C;
        15'h3AFE: data = 12'h75C;
        15'h3AFF: data = 12'h747;
        15'h3B00: data = 12'h73C;
        15'h3B01: data = 12'h729;
        15'h3B02: data = 12'h726;
        15'h3B03: data = 12'h71C;
        15'h3B04: data = 12'h711;
        15'h3B05: data = 12'h709;
        15'h3B06: data = 12'h6FC;
        15'h3B07: data = 12'h6EA;
        15'h3B08: data = 12'h6DA;
        15'h3B09: data = 12'h6C5;
        15'h3B0A: data = 12'h6B3;
        15'h3B0B: data = 12'h6A6;
        15'h3B0C: data = 12'h696;
        15'h3B0D: data = 12'h68B;
        15'h3B0E: data = 12'h682;
        15'h3B0F: data = 12'h677;
        15'h3B10: data = 12'h66A;
        15'h3B11: data = 12'h65B;
        15'h3B12: data = 12'h647;
        15'h3B13: data = 12'h634;
        15'h3B14: data = 12'h625;
        15'h3B15: data = 12'h60A;
        15'h3B16: data = 12'h5F6;
        15'h3B17: data = 12'h5E4;
        15'h3B18: data = 12'h5CF;
        15'h3B19: data = 12'h5BE;
        15'h3B1A: data = 12'h5B6;
        15'h3B1B: data = 12'h5A4;
        15'h3B1C: data = 12'h597;
        15'h3B1D: data = 12'h584;
        15'h3B1E: data = 12'h574;
        15'h3B1F: data = 12'h567;
        15'h3B20: data = 12'h556;
        15'h3B21: data = 12'h542;
        15'h3B22: data = 12'h52B;
        15'h3B23: data = 12'h518;
        15'h3B24: data = 12'h504;
        15'h3B25: data = 12'h4F1;
        15'h3B26: data = 12'h4D7;
        15'h3B27: data = 12'h4BA;
        15'h3B28: data = 12'h4AC;
        15'h3B29: data = 12'h492;
        15'h3B2A: data = 12'h47A;
        15'h3B2B: data = 12'h463;
        15'h3B2C: data = 12'h451;
        15'h3B2D: data = 12'h43D;
        15'h3B2E: data = 12'h42C;
        15'h3B2F: data = 12'h419;
        15'h3B30: data = 12'h402;
        15'h3B31: data = 12'h3E9;
        15'h3B32: data = 12'h3D7;
        15'h3B33: data = 12'h3C3;
        15'h3B34: data = 12'h3B1;
        15'h3B35: data = 12'h398;
        15'h3B36: data = 12'h387;
        15'h3B37: data = 12'h371;
        15'h3B38: data = 12'h35D;
        15'h3B39: data = 12'h348;
        15'h3B3A: data = 12'h330;
        15'h3B3B: data = 12'h31C;
        15'h3B3C: data = 12'h301;
        15'h3B3D: data = 12'h2EE;
        15'h3B3E: data = 12'h2DA;
        15'h3B3F: data = 12'h2C7;
        15'h3B40: data = 12'h2AB;
        15'h3B41: data = 12'h292;
        15'h3B42: data = 12'h27E;
        15'h3B43: data = 12'h264;
        15'h3B44: data = 12'h24B;
        15'h3B45: data = 12'h234;
        15'h3B46: data = 12'h21D;
        15'h3B47: data = 12'h205;
        15'h3B48: data = 12'h1F0;
        15'h3B49: data = 12'h1D8;
        15'h3B4A: data = 12'h1C0;
        15'h3B4B: data = 12'h1AC;
        15'h3B4C: data = 12'h193;
        15'h3B4D: data = 12'h17C;
        15'h3B4E: data = 12'h166;
        15'h3B4F: data = 12'h14E;
        15'h3B50: data = 12'h137;
        15'h3B51: data = 12'h11B;
        15'h3B52: data = 12'h107;
        15'h3B53: data = 12'h0F5;
        15'h3B54: data = 12'h0D9;
        15'h3B55: data = 12'h0BF;
        15'h3B56: data = 12'h0A6;
        15'h3B57: data = 12'h093;
        15'h3B58: data = 12'h07C;
        15'h3B59: data = 12'h062;
        15'h3B5A: data = 12'h04E;
        15'h3B5B: data = 12'h680;
        15'h3B5C: data = 12'h7CF;
        15'h3B5D: data = 12'h7BA;
        15'h3B5E: data = 12'h7A5;
        15'h3B5F: data = 12'h78C;
        15'h3B60: data = 12'h776;
        15'h3B61: data = 12'h75A;
        15'h3B62: data = 12'h74A;
        15'h3B63: data = 12'h734;
        15'h3B64: data = 12'h71E;
        15'h3B65: data = 12'h708;
        15'h3B66: data = 12'h6EB;
        15'h3B67: data = 12'h6D9;
        15'h3B68: data = 12'h6C2;
        15'h3B69: data = 12'h6AA;
        15'h3B6A: data = 12'h68F;
        15'h3B6B: data = 12'h67B;
        15'h3B6C: data = 12'h664;
        15'h3B6D: data = 12'h654;
        15'h3B6E: data = 12'h63A;
        15'h3B6F: data = 12'h624;
        15'h3B70: data = 12'h60F;
        15'h3B71: data = 12'h5F7;
        15'h3B72: data = 12'h5DF;
        15'h3B73: data = 12'h5C9;
        15'h3B74: data = 12'h5B3;
        15'h3B75: data = 12'h59B;
        15'h3B76: data = 12'h581;
        15'h3B77: data = 12'h56C;
        15'h3B78: data = 12'h55D;
        15'h3B79: data = 12'h544;
        15'h3B7A: data = 12'h531;
        15'h3B7B: data = 12'h51B;
        15'h3B7C: data = 12'h507;
        15'h3B7D: data = 12'h4F4;
        15'h3B7E: data = 12'h4DD;
        15'h3B7F: data = 12'h4C9;
        15'h3B80: data = 12'h4B7;
        15'h3B81: data = 12'h4A4;
        15'h3B82: data = 12'h492;
        15'h3B83: data = 12'h47F;
        15'h3B84: data = 12'h46C;
        15'h3B85: data = 12'h45E;
        15'h3B86: data = 12'h44D;
        15'h3B87: data = 12'h43A;
        15'h3B88: data = 12'h42C;
        15'h3B89: data = 12'h418;
        15'h3B8A: data = 12'h407;
        15'h3B8B: data = 12'h3F7;
        15'h3B8C: data = 12'h3EC;
        15'h3B8D: data = 12'h3D2;
        15'h3B8E: data = 12'h3C0;
        15'h3B8F: data = 12'h3AC;
        15'h3B90: data = 12'h396;
        15'h3B91: data = 12'h38D;
        15'h3B92: data = 12'h376;
        15'h3B93: data = 12'h363;
        15'h3B94: data = 12'h34F;
        15'h3B95: data = 12'h33E;
        15'h3B96: data = 12'h32E;
        15'h3B97: data = 12'h31C;
        15'h3B98: data = 12'h310;
        15'h3B99: data = 12'h2FE;
        15'h3B9A: data = 12'h2F3;
        15'h3B9B: data = 12'h2E7;
        15'h3B9C: data = 12'h2D8;
        15'h3B9D: data = 12'h2D8;
        15'h3B9E: data = 12'h2C7;
        15'h3B9F: data = 12'h2BB;
        15'h3BA0: data = 12'h2AA;
        15'h3BA1: data = 12'h2A0;
        15'h3BA2: data = 12'h297;
        15'h3BA3: data = 12'h284;
        15'h3BA4: data = 12'h27B;
        15'h3BA5: data = 12'h26B;
        15'h3BA6: data = 12'h25C;
        15'h3BA7: data = 12'h24B;
        15'h3BA8: data = 12'h23C;
        15'h3BA9: data = 12'h22C;
        15'h3BAA: data = 12'h220;
        15'h3BAB: data = 12'h214;
        15'h3BAC: data = 12'h213;
        15'h3BAD: data = 12'h20B;
        15'h3BAE: data = 12'h207;
        15'h3BAF: data = 12'h1FD;
        15'h3BB0: data = 12'h1F7;
        15'h3BB1: data = 12'h1F1;
        15'h3BB2: data = 12'h1EC;
        15'h3BB3: data = 12'h1DF;
        15'h3BB4: data = 12'h1D4;
        15'h3BB5: data = 12'h1C7;
        15'h3BB6: data = 12'h1BB;
        15'h3BB7: data = 12'h1B7;
        15'h3BB8: data = 12'h1AB;
        15'h3BB9: data = 12'h1A3;
        15'h3BBA: data = 12'h199;
        15'h3BBB: data = 12'h195;
        15'h3BBC: data = 12'h194;
        15'h3BBD: data = 12'h18F;
        15'h3BBE: data = 12'h18F;
        15'h3BBF: data = 12'h18A;
        15'h3BC0: data = 12'h18C;
        15'h3BC1: data = 12'h188;
        15'h3BC2: data = 12'h188;
        15'h3BC3: data = 12'h17F;
        15'h3BC4: data = 12'h17D;
        15'h3BC5: data = 12'h174;
        15'h3BC6: data = 12'h16E;
        15'h3BC7: data = 12'h16A;
        15'h3BC8: data = 12'h160;
        15'h3BC9: data = 12'h161;
        15'h3BCA: data = 12'h15E;
        15'h3BCB: data = 12'h15F;
        15'h3BCC: data = 12'h155;
        15'h3BCD: data = 12'h15C;
        15'h3BCE: data = 12'h15E;
        15'h3BCF: data = 12'h164;
        15'h3BD0: data = 12'h168;
        15'h3BD1: data = 12'h168;
        15'h3BD2: data = 12'h168;
        15'h3BD3: data = 12'h170;
        15'h3BD4: data = 12'h16E;
        15'h3BD5: data = 12'h16C;
        15'h3BD6: data = 12'h16A;
        15'h3BD7: data = 12'h162;
        15'h3BD8: data = 12'h168;
        15'h3BD9: data = 12'h165;
        15'h3BDA: data = 12'h16C;
        15'h3BDB: data = 12'h16F;
        15'h3BDC: data = 12'h171;
        15'h3BDD: data = 12'h17A;
        15'h3BDE: data = 12'h184;
        15'h3BDF: data = 12'h187;
        15'h3BE0: data = 12'h194;
        15'h3BE1: data = 12'h197;
        15'h3BE2: data = 12'h1A0;
        15'h3BE3: data = 12'h1A2;
        15'h3BE4: data = 12'h1AC;
        15'h3BE5: data = 12'h1B1;
        15'h3BE6: data = 12'h1B2;
        15'h3BE7: data = 12'h1B4;
        15'h3BE8: data = 12'h1B5;
        15'h3BE9: data = 12'h1B9;
        15'h3BEA: data = 12'h1C0;
        15'h3BEB: data = 12'h1C9;
        15'h3BEC: data = 12'h1D2;
        15'h3BED: data = 12'h1DB;
        15'h3BEE: data = 12'h1E7;
        15'h3BEF: data = 12'h1F9;
        15'h3BF0: data = 12'h201;
        15'h3BF1: data = 12'h20F;
        15'h3BF2: data = 12'h21F;
        15'h3BF3: data = 12'h220;
        15'h3BF4: data = 12'h234;
        15'h3BF5: data = 12'h238;
        15'h3BF6: data = 12'h247;
        15'h3BF7: data = 12'h24D;
        15'h3BF8: data = 12'h258;
        15'h3BF9: data = 12'h25D;
        15'h3BFA: data = 12'h266;
        15'h3BFB: data = 12'h269;
        15'h3BFC: data = 12'h279;
        15'h3BFD: data = 12'h289;
        15'h3BFE: data = 12'h291;
        15'h3BFF: data = 12'h2A3;
        15'h3C00: data = 12'h2B1;
        15'h3C01: data = 12'h2C7;
        15'h3C02: data = 12'h2D8;
        15'h3C03: data = 12'h2E6;
        15'h3C04: data = 12'h2F6;
        15'h3C05: data = 12'h308;
        15'h3C06: data = 12'h31A;
        15'h3C07: data = 12'h327;
        15'h3C08: data = 12'h339;
        15'h3C09: data = 12'h347;
        15'h3C0A: data = 12'h355;
        15'h3C0B: data = 12'h360;
        15'h3C0C: data = 12'h36E;
        15'h3C0D: data = 12'h379;
        15'h3C0E: data = 12'h38D;
        15'h3C0F: data = 12'h394;
        15'h3C10: data = 12'h3AB;
        15'h3C11: data = 12'h3B7;
        15'h3C12: data = 12'h3C7;
        15'h3C13: data = 12'h3DE;
        15'h3C14: data = 12'h3F1;
        15'h3C15: data = 12'h404;
        15'h3C16: data = 12'h41F;
        15'h3C17: data = 12'h431;
        15'h3C18: data = 12'h44A;
        15'h3C19: data = 12'h45E;
        15'h3C1A: data = 12'h46F;
        15'h3C1B: data = 12'h484;
        15'h3C1C: data = 12'h497;
        15'h3C1D: data = 12'h4AB;
        15'h3C1E: data = 12'h4B7;
        15'h3C1F: data = 12'h4CB;
        15'h3C20: data = 12'h4E3;
        15'h3C21: data = 12'h4F2;
        15'h3C22: data = 12'h506;
        15'h3C23: data = 12'h513;
        15'h3C24: data = 12'h524;
        15'h3C25: data = 12'h53B;
        15'h3C26: data = 12'h553;
        15'h3C27: data = 12'h565;
        15'h3C28: data = 12'h578;
        15'h3C29: data = 12'h58D;
        15'h3C2A: data = 12'h5A5;
        15'h3C2B: data = 12'h5BC;
        15'h3C2C: data = 12'h5D1;
        15'h3C2D: data = 12'h5EE;
        15'h3C2E: data = 12'h607;
        15'h3C2F: data = 12'h61F;
        15'h3C30: data = 12'h636;
        15'h3C31: data = 12'h64E;
        15'h3C32: data = 12'h663;
        15'h3C33: data = 12'h677;
        15'h3C34: data = 12'h692;
        15'h3C35: data = 12'h6A3;
        15'h3C36: data = 12'h6B6;
        15'h3C37: data = 12'h6D2;
        15'h3C38: data = 12'h6DF;
        15'h3C39: data = 12'h6F3;
        15'h3C3A: data = 12'h703;
        15'h3C3B: data = 12'h71E;
        15'h3C3C: data = 12'h737;
        15'h3C3D: data = 12'h744;
        15'h3C3E: data = 12'h75C;
        15'h3C3F: data = 12'h776;
        15'h3C40: data = 12'h794;
        15'h3C41: data = 12'h7A3;
        15'h3C42: data = 12'h7C0;
        15'h3C43: data = 12'h7DC;
        15'h3C44: data = 12'h7F1;
        15'h3C45: data = 12'h806;
        15'h3C46: data = 12'h078;
        15'h3C47: data = 12'h092;
        15'h3C48: data = 12'h0A6;
        15'h3C49: data = 12'h0BC;
        15'h3C4A: data = 12'h0D1;
        15'h3C4B: data = 12'h0EB;
        15'h3C4C: data = 12'h0FF;
        15'h3C4D: data = 12'h112;
        15'h3C4E: data = 12'h127;
        15'h3C4F: data = 12'h141;
        15'h3C50: data = 12'h155;
        15'h3C51: data = 12'h165;
        15'h3C52: data = 12'h17C;
        15'h3C53: data = 12'h196;
        15'h3C54: data = 12'h1AB;
        15'h3C55: data = 12'h1BD;
        15'h3C56: data = 12'h1D7;
        15'h3C57: data = 12'h1EC;
        15'h3C58: data = 12'h205;
        15'h3C59: data = 12'h21B;
        15'h3C5A: data = 12'h231;
        15'h3C5B: data = 12'h249;
        15'h3C5C: data = 12'h265;
        15'h3C5D: data = 12'h27B;
        15'h3C5E: data = 12'h28E;
        15'h3C5F: data = 12'h2AE;
        15'h3C60: data = 12'h2C6;
        15'h3C61: data = 12'h2DC;
        15'h3C62: data = 12'h2FB;
        15'h3C63: data = 12'h30E;
        15'h3C64: data = 12'h32B;
        15'h3C65: data = 12'h33D;
        15'h3C66: data = 12'h351;
        15'h3C67: data = 12'h36C;
        15'h3C68: data = 12'h37F;
        15'h3C69: data = 12'h39B;
        15'h3C6A: data = 12'h3AD;
        15'h3C6B: data = 12'h3C4;
        15'h3C6C: data = 12'h3D6;
        15'h3C6D: data = 12'h3EF;
        15'h3C6E: data = 12'h3FE;
        15'h3C6F: data = 12'h414;
        15'h3C70: data = 12'h42B;
        15'h3C71: data = 12'h442;
        15'h3C72: data = 12'h44E;
        15'h3C73: data = 12'h461;
        15'h3C74: data = 12'h477;
        15'h3C75: data = 12'h48F;
        15'h3C76: data = 12'h4A3;
        15'h3C77: data = 12'h4B1;
        15'h3C78: data = 12'h4C1;
        15'h3C79: data = 12'h4D6;
        15'h3C7A: data = 12'h4EA;
        15'h3C7B: data = 12'h505;
        15'h3C7C: data = 12'h513;
        15'h3C7D: data = 12'h524;
        15'h3C7E: data = 12'h53A;
        15'h3C7F: data = 12'h549;
        15'h3C80: data = 12'h55A;
        15'h3C81: data = 12'h56D;
        15'h3C82: data = 12'h585;
        15'h3C83: data = 12'h593;
        15'h3C84: data = 12'h5AA;
        15'h3C85: data = 12'h5BA;
        15'h3C86: data = 12'h5CA;
        15'h3C87: data = 12'h5DA;
        15'h3C88: data = 12'h5F3;
        15'h3C89: data = 12'h600;
        15'h3C8A: data = 12'h613;
        15'h3C8B: data = 12'h623;
        15'h3C8C: data = 12'h634;
        15'h3C8D: data = 12'h645;
        15'h3C8E: data = 12'h659;
        15'h3C8F: data = 12'h66D;
        15'h3C90: data = 12'h67B;
        15'h3C91: data = 12'h689;
        15'h3C92: data = 12'h69A;
        15'h3C93: data = 12'h6AD;
        15'h3C94: data = 12'h6BB;
        15'h3C95: data = 12'h6CA;
        15'h3C96: data = 12'h6D8;
        15'h3C97: data = 12'h6DE;
        15'h3C98: data = 12'h6F0;
        15'h3C99: data = 12'h6FF;
        15'h3C9A: data = 12'h70A;
        15'h3C9B: data = 12'h716;
        15'h3C9C: data = 12'h723;
        15'h3C9D: data = 12'h738;
        15'h3C9E: data = 12'h73B;
        15'h3C9F: data = 12'h74A;
        15'h3CA0: data = 12'h74F;
        15'h3CA1: data = 12'h75F;
        15'h3CA2: data = 12'h766;
        15'h3CA3: data = 12'h777;
        15'h3CA4: data = 12'h77F;
        15'h3CA5: data = 12'h78C;
        15'h3CA6: data = 12'h792;
        15'h3CA7: data = 12'h79C;
        15'h3CA8: data = 12'h7A3;
        15'h3CA9: data = 12'h7AE;
        15'h3CAA: data = 12'h7B5;
        15'h3CAB: data = 12'h7BE;
        15'h3CAC: data = 12'h7C1;
        15'h3CAD: data = 12'h7C7;
        15'h3CAE: data = 12'h7CE;
        15'h3CAF: data = 12'h7D7;
        15'h3CB0: data = 12'h7DF;
        15'h3CB1: data = 12'h7E6;
        15'h3CB2: data = 12'h7E9;
        15'h3CB3: data = 12'h7F3;
        15'h3CB4: data = 12'h7F9;
        15'h3CB5: data = 12'h7FC;
        15'h3CB6: data = 12'h7FF;
        15'h3CB7: data = 12'h805;
        15'h3CB8: data = 12'h74D;
        15'h3CB9: data = 12'h087;
        15'h3CBA: data = 12'h08D;
        15'h3CBB: data = 12'h095;
        15'h3CBC: data = 12'h094;
        15'h3CBD: data = 12'h09F;
        15'h3CBE: data = 12'h0A1;
        15'h3CBF: data = 12'h0AA;
        15'h3CC0: data = 12'h0AD;
        15'h3CC1: data = 12'h0AD;
        15'h3CC2: data = 12'h0B5;
        15'h3CC3: data = 12'h0B9;
        15'h3CC4: data = 12'h0BD;
        15'h3CC5: data = 12'h0BE;
        15'h3CC6: data = 12'h0CA;
        15'h3CC7: data = 12'h0CF;
        15'h3CC8: data = 12'h0CF;
        15'h3CC9: data = 12'h0D1;
        15'h3CCA: data = 12'h0D1;
        15'h3CCB: data = 12'h0D6;
        15'h3CCC: data = 12'h0D5;
        15'h3CCD: data = 12'h0CB;
        15'h3CCE: data = 12'h0C8;
        15'h3CCF: data = 12'h0CA;
        15'h3CD0: data = 12'h0C8;
        15'h3CD1: data = 12'h0BC;
        15'h3CD2: data = 12'h0B5;
        15'h3CD3: data = 12'h0B4;
        15'h3CD4: data = 12'h0AD;
        15'h3CD5: data = 12'h0AD;
        15'h3CD6: data = 12'h0AA;
        15'h3CD7: data = 12'h0AD;
        15'h3CD8: data = 12'h0AE;
        15'h3CD9: data = 12'h0B4;
        15'h3CDA: data = 12'h0AC;
        15'h3CDB: data = 12'h0A5;
        15'h3CDC: data = 12'h0A3;
        15'h3CDD: data = 12'h098;
        15'h3CDE: data = 12'h08B;
        15'h3CDF: data = 12'h07E;
        15'h3CE0: data = 12'h075;
        15'h3CE1: data = 12'h075;
        15'h3CE2: data = 12'h070;
        15'h3CE3: data = 12'h06F;
        15'h3CE4: data = 12'h070;
        15'h3CE5: data = 12'h06A;
        15'h3CE6: data = 12'h05F;
        15'h3CE7: data = 12'h057;
        15'h3CE8: data = 12'h044;
        15'h3CE9: data = 12'h7BC;
        15'h3CEA: data = 12'h7AE;
        15'h3CEB: data = 12'h7A5;
        15'h3CEC: data = 12'h7A2;
        15'h3CED: data = 12'h798;
        15'h3CEE: data = 12'h794;
        15'h3CEF: data = 12'h78B;
        15'h3CF0: data = 12'h779;
        15'h3CF1: data = 12'h76A;
        15'h3CF2: data = 12'h758;
        15'h3CF3: data = 12'h741;
        15'h3CF4: data = 12'h735;
        15'h3CF5: data = 12'h72C;
        15'h3CF6: data = 12'h727;
        15'h3CF7: data = 12'h71C;
        15'h3CF8: data = 12'h710;
        15'h3CF9: data = 12'h70C;
        15'h3CFA: data = 12'h6FC;
        15'h3CFB: data = 12'h6EC;
        15'h3CFC: data = 12'h6D9;
        15'h3CFD: data = 12'h6C6;
        15'h3CFE: data = 12'h6B0;
        15'h3CFF: data = 12'h6A3;
        15'h3D00: data = 12'h694;
        15'h3D01: data = 12'h68B;
        15'h3D02: data = 12'h67F;
        15'h3D03: data = 12'h674;
        15'h3D04: data = 12'h669;
        15'h3D05: data = 12'h655;
        15'h3D06: data = 12'h646;
        15'h3D07: data = 12'h632;
        15'h3D08: data = 12'h629;
        15'h3D09: data = 12'h60E;
        15'h3D0A: data = 12'h5F9;
        15'h3D0B: data = 12'h5E5;
        15'h3D0C: data = 12'h5CF;
        15'h3D0D: data = 12'h5BD;
        15'h3D0E: data = 12'h5B1;
        15'h3D0F: data = 12'h5A0;
        15'h3D10: data = 12'h592;
        15'h3D11: data = 12'h57F;
        15'h3D12: data = 12'h571;
        15'h3D13: data = 12'h566;
        15'h3D14: data = 12'h552;
        15'h3D15: data = 12'h541;
        15'h3D16: data = 12'h52C;
        15'h3D17: data = 12'h516;
        15'h3D18: data = 12'h506;
        15'h3D19: data = 12'h4F3;
        15'h3D1A: data = 12'h4D9;
        15'h3D1B: data = 12'h4C1;
        15'h3D1C: data = 12'h4AC;
        15'h3D1D: data = 12'h492;
        15'h3D1E: data = 12'h47C;
        15'h3D1F: data = 12'h465;
        15'h3D20: data = 12'h452;
        15'h3D21: data = 12'h43C;
        15'h3D22: data = 12'h42A;
        15'h3D23: data = 12'h413;
        15'h3D24: data = 12'h3FF;
        15'h3D25: data = 12'h3E6;
        15'h3D26: data = 12'h3D0;
        15'h3D27: data = 12'h3BF;
        15'h3D28: data = 12'h3AB;
        15'h3D29: data = 12'h392;
        15'h3D2A: data = 12'h380;
        15'h3D2B: data = 12'h36A;
        15'h3D2C: data = 12'h356;
        15'h3D2D: data = 12'h33F;
        15'h3D2E: data = 12'h329;
        15'h3D2F: data = 12'h317;
        15'h3D30: data = 12'h300;
        15'h3D31: data = 12'h2EC;
        15'h3D32: data = 12'h2D5;
        15'h3D33: data = 12'h2C1;
        15'h3D34: data = 12'h2A5;
        15'h3D35: data = 12'h28E;
        15'h3D36: data = 12'h27E;
        15'h3D37: data = 12'h264;
        15'h3D38: data = 12'h24B;
        15'h3D39: data = 12'h234;
        15'h3D3A: data = 12'h21D;
        15'h3D3B: data = 12'h205;
        15'h3D3C: data = 12'h1F1;
        15'h3D3D: data = 12'h1D6;
        15'h3D3E: data = 12'h1C2;
        15'h3D3F: data = 12'h1AA;
        15'h3D40: data = 12'h193;
        15'h3D41: data = 12'h17C;
        15'h3D42: data = 12'h165;
        15'h3D43: data = 12'h14E;
        15'h3D44: data = 12'h139;
        15'h3D45: data = 12'h11C;
        15'h3D46: data = 12'h107;
        15'h3D47: data = 12'h0F5;
        15'h3D48: data = 12'h0D6;
        15'h3D49: data = 12'h0C1;
        15'h3D4A: data = 12'h0A7;
        15'h3D4B: data = 12'h08E;
        15'h3D4C: data = 12'h07D;
        15'h3D4D: data = 12'h065;
        15'h3D4E: data = 12'h04E;
        15'h3D4F: data = 12'h7E0;
        15'h3D50: data = 12'h7CD;
        15'h3D51: data = 12'h7BB;
        15'h3D52: data = 12'h7A4;
        15'h3D53: data = 12'h78D;
        15'h3D54: data = 12'h773;
        15'h3D55: data = 12'h758;
        15'h3D56: data = 12'h748;
        15'h3D57: data = 12'h736;
        15'h3D58: data = 12'h71C;
        15'h3D59: data = 12'h704;
        15'h3D5A: data = 12'h6E9;
        15'h3D5B: data = 12'h6D9;
        15'h3D5C: data = 12'h6C1;
        15'h3D5D: data = 12'h6AB;
        15'h3D5E: data = 12'h695;
        15'h3D5F: data = 12'h67E;
        15'h3D60: data = 12'h666;
        15'h3D61: data = 12'h64F;
        15'h3D62: data = 12'h63C;
        15'h3D63: data = 12'h62A;
        15'h3D64: data = 12'h611;
        15'h3D65: data = 12'h5F5;
        15'h3D66: data = 12'h5DF;
        15'h3D67: data = 12'h5CB;
        15'h3D68: data = 12'h5B4;
        15'h3D69: data = 12'h59A;
        15'h3D6A: data = 12'h582;
        15'h3D6B: data = 12'h56F;
        15'h3D6C: data = 12'h55A;
        15'h3D6D: data = 12'h546;
        15'h3D6E: data = 12'h530;
        15'h3D6F: data = 12'h51C;
        15'h3D70: data = 12'h505;
        15'h3D71: data = 12'h4F3;
        15'h3D72: data = 12'h4E0;
        15'h3D73: data = 12'h4CA;
        15'h3D74: data = 12'h4B5;
        15'h3D75: data = 12'h4A0;
        15'h3D76: data = 12'h492;
        15'h3D77: data = 12'h47D;
        15'h3D78: data = 12'h469;
        15'h3D79: data = 12'h459;
        15'h3D7A: data = 12'h44E;
        15'h3D7B: data = 12'h43C;
        15'h3D7C: data = 12'h42E;
        15'h3D7D: data = 12'h418;
        15'h3D7E: data = 12'h406;
        15'h3D7F: data = 12'h3F9;
        15'h3D80: data = 12'h3EA;
        15'h3D81: data = 12'h3D0;
        15'h3D82: data = 12'h3C2;
        15'h3D83: data = 12'h3AC;
        15'h3D84: data = 12'h399;
        15'h3D85: data = 12'h390;
        15'h3D86: data = 12'h375;
        15'h3D87: data = 12'h362;
        15'h3D88: data = 12'h34D;
        15'h3D89: data = 12'h33E;
        15'h3D8A: data = 12'h32D;
        15'h3D8B: data = 12'h31D;
        15'h3D8C: data = 12'h30D;
        15'h3D8D: data = 12'h2FD;
        15'h3D8E: data = 12'h2F2;
        15'h3D8F: data = 12'h2E4;
        15'h3D90: data = 12'h2DA;
        15'h3D91: data = 12'h2D5;
        15'h3D92: data = 12'h2C6;
        15'h3D93: data = 12'h2BC;
        15'h3D94: data = 12'h2AB;
        15'h3D95: data = 12'h29C;
        15'h3D96: data = 12'h293;
        15'h3D97: data = 12'h282;
        15'h3D98: data = 12'h279;
        15'h3D99: data = 12'h266;
        15'h3D9A: data = 12'h25A;
        15'h3D9B: data = 12'h248;
        15'h3D9C: data = 12'h238;
        15'h3D9D: data = 12'h22A;
        15'h3D9E: data = 12'h220;
        15'h3D9F: data = 12'h217;
        15'h3DA0: data = 12'h20F;
        15'h3DA1: data = 12'h20D;
        15'h3DA2: data = 12'h209;
        15'h3DA3: data = 12'h1FE;
        15'h3DA4: data = 12'h1F9;
        15'h3DA5: data = 12'h1F4;
        15'h3DA6: data = 12'h1EC;
        15'h3DA7: data = 12'h1DE;
        15'h3DA8: data = 12'h1D0;
        15'h3DA9: data = 12'h1C8;
        15'h3DAA: data = 12'h1BB;
        15'h3DAB: data = 12'h1B3;
        15'h3DAC: data = 12'h1A9;
        15'h3DAD: data = 12'h19F;
        15'h3DAE: data = 12'h19A;
        15'h3DAF: data = 12'h192;
        15'h3DB0: data = 12'h195;
        15'h3DB1: data = 12'h193;
        15'h3DB2: data = 12'h18C;
        15'h3DB3: data = 12'h18A;
        15'h3DB4: data = 12'h18C;
        15'h3DB5: data = 12'h187;
        15'h3DB6: data = 12'h188;
        15'h3DB7: data = 12'h181;
        15'h3DB8: data = 12'h17E;
        15'h3DB9: data = 12'h172;
        15'h3DBA: data = 12'h16F;
        15'h3DBB: data = 12'h169;
        15'h3DBC: data = 12'h161;
        15'h3DBD: data = 12'h15C;
        15'h3DBE: data = 12'h15D;
        15'h3DBF: data = 12'h15E;
        15'h3DC0: data = 12'h158;
        15'h3DC1: data = 12'h15D;
        15'h3DC2: data = 12'h15F;
        15'h3DC3: data = 12'h164;
        15'h3DC4: data = 12'h164;
        15'h3DC5: data = 12'h169;
        15'h3DC6: data = 12'h16A;
        15'h3DC7: data = 12'h16F;
        15'h3DC8: data = 12'h170;
        15'h3DC9: data = 12'h16D;
        15'h3DCA: data = 12'h168;
        15'h3DCB: data = 12'h163;
        15'h3DCC: data = 12'h167;
        15'h3DCD: data = 12'h164;
        15'h3DCE: data = 12'h16D;
        15'h3DCF: data = 12'h16D;
        15'h3DD0: data = 12'h16D;
        15'h3DD1: data = 12'h17C;
        15'h3DD2: data = 12'h185;
        15'h3DD3: data = 12'h189;
        15'h3DD4: data = 12'h193;
        15'h3DD5: data = 12'h197;
        15'h3DD6: data = 12'h19F;
        15'h3DD7: data = 12'h1A2;
        15'h3DD8: data = 12'h1AC;
        15'h3DD9: data = 12'h1B3;
        15'h3DDA: data = 12'h1B2;
        15'h3DDB: data = 12'h1B3;
        15'h3DDC: data = 12'h1B9;
        15'h3DDD: data = 12'h1BC;
        15'h3DDE: data = 12'h1BF;
        15'h3DDF: data = 12'h1C6;
        15'h3DE0: data = 12'h1CE;
        15'h3DE1: data = 12'h1D8;
        15'h3DE2: data = 12'h1E8;
        15'h3DE3: data = 12'h1F6;
        15'h3DE4: data = 12'h200;
        15'h3DE5: data = 12'h20D;
        15'h3DE6: data = 12'h223;
        15'h3DE7: data = 12'h220;
        15'h3DE8: data = 12'h22F;
        15'h3DE9: data = 12'h239;
        15'h3DEA: data = 12'h246;
        15'h3DEB: data = 12'h24C;
        15'h3DEC: data = 12'h259;
        15'h3DED: data = 12'h260;
        15'h3DEE: data = 12'h26A;
        15'h3DEF: data = 12'h26B;
        15'h3DF0: data = 12'h27B;
        15'h3DF1: data = 12'h289;
        15'h3DF2: data = 12'h292;
        15'h3DF3: data = 12'h2A4;
        15'h3DF4: data = 12'h2B8;
        15'h3DF5: data = 12'h2C7;
        15'h3DF6: data = 12'h2DA;
        15'h3DF7: data = 12'h2E3;
        15'h3DF8: data = 12'h2F9;
        15'h3DF9: data = 12'h309;
        15'h3DFA: data = 12'h318;
        15'h3DFB: data = 12'h324;
        15'h3DFC: data = 12'h337;
        15'h3DFD: data = 12'h345;
        15'h3DFE: data = 12'h350;
        15'h3DFF: data = 12'h362;
        15'h3E00: data = 12'h36E;
        15'h3E01: data = 12'h378;
        15'h3E02: data = 12'h38C;
        15'h3E03: data = 12'h394;
        15'h3E04: data = 12'h3A5;
        15'h3E05: data = 12'h3B4;
        15'h3E06: data = 12'h3C6;
        15'h3E07: data = 12'h3DE;
        15'h3E08: data = 12'h3EF;
        15'h3E09: data = 12'h402;
        15'h3E0A: data = 12'h41B;
        15'h3E0B: data = 12'h431;
        15'h3E0C: data = 12'h447;
        15'h3E0D: data = 12'h459;
        15'h3E0E: data = 12'h46D;
        15'h3E0F: data = 12'h481;
        15'h3E10: data = 12'h495;
        15'h3E11: data = 12'h4A8;
        15'h3E12: data = 12'h4B8;
        15'h3E13: data = 12'h4CE;
        15'h3E14: data = 12'h4E2;
        15'h3E15: data = 12'h4F4;
        15'h3E16: data = 12'h508;
        15'h3E17: data = 12'h51A;
        15'h3E18: data = 12'h524;
        15'h3E19: data = 12'h53B;
        15'h3E1A: data = 12'h54D;
        15'h3E1B: data = 12'h564;
        15'h3E1C: data = 12'h575;
        15'h3E1D: data = 12'h58C;
        15'h3E1E: data = 12'h5A3;
        15'h3E1F: data = 12'h5BC;
        15'h3E20: data = 12'h5D0;
        15'h3E21: data = 12'h5E8;
        15'h3E22: data = 12'h605;
        15'h3E23: data = 12'h61C;
        15'h3E24: data = 12'h636;
        15'h3E25: data = 12'h649;
        15'h3E26: data = 12'h666;
        15'h3E27: data = 12'h678;
        15'h3E28: data = 12'h691;
        15'h3E29: data = 12'h6A1;
        15'h3E2A: data = 12'h6B6;
        15'h3E2B: data = 12'h6D0;
        15'h3E2C: data = 12'h6DD;
        15'h3E2D: data = 12'h6F4;
        15'h3E2E: data = 12'h706;
        15'h3E2F: data = 12'h71C;
        15'h3E30: data = 12'h734;
        15'h3E31: data = 12'h742;
        15'h3E32: data = 12'h75B;
        15'h3E33: data = 12'h774;
        15'h3E34: data = 12'h790;
        15'h3E35: data = 12'h7A1;
        15'h3E36: data = 12'h7BE;
        15'h3E37: data = 12'h7DD;
        15'h3E38: data = 12'h7F2;
        15'h3E39: data = 12'h807;
        15'h3E3A: data = 12'h077;
        15'h3E3B: data = 12'h08D;
        15'h3E3C: data = 12'h0A2;
        15'h3E3D: data = 12'h0BC;
        15'h3E3E: data = 12'h0D6;
        15'h3E3F: data = 12'h0EA;
        15'h3E40: data = 12'h101;
        15'h3E41: data = 12'h113;
        15'h3E42: data = 12'h129;
        15'h3E43: data = 12'h144;
        15'h3E44: data = 12'h155;
        15'h3E45: data = 12'h168;
        15'h3E46: data = 12'h17B;
        15'h3E47: data = 12'h196;
        15'h3E48: data = 12'h1AC;
        15'h3E49: data = 12'h1BB;
        15'h3E4A: data = 12'h1D7;
        15'h3E4B: data = 12'h1EB;
        15'h3E4C: data = 12'h205;
        15'h3E4D: data = 12'h217;
        15'h3E4E: data = 12'h230;
        15'h3E4F: data = 12'h24B;
        15'h3E50: data = 12'h261;
        15'h3E51: data = 12'h279;
        15'h3E52: data = 12'h290;
        15'h3E53: data = 12'h2AB;
        15'h3E54: data = 12'h2C3;
        15'h3E55: data = 12'h2DE;
        15'h3E56: data = 12'h2F8;
        15'h3E57: data = 12'h30E;
        15'h3E58: data = 12'h328;
        15'h3E59: data = 12'h339;
        15'h3E5A: data = 12'h34F;
        15'h3E5B: data = 12'h36B;
        15'h3E5C: data = 12'h37F;
        15'h3E5D: data = 12'h39A;
        15'h3E5E: data = 12'h3AA;
        15'h3E5F: data = 12'h3C0;
        15'h3E60: data = 12'h3D5;
        15'h3E61: data = 12'h3F2;
        15'h3E62: data = 12'h3FE;
        15'h3E63: data = 12'h414;
        15'h3E64: data = 12'h42E;
        15'h3E65: data = 12'h442;
        15'h3E66: data = 12'h451;
        15'h3E67: data = 12'h462;
        15'h3E68: data = 12'h479;
        15'h3E69: data = 12'h490;
        15'h3E6A: data = 12'h4A2;
        15'h3E6B: data = 12'h4B3;
        15'h3E6C: data = 12'h4C1;
        15'h3E6D: data = 12'h4D5;
        15'h3E6E: data = 12'h4EA;
        15'h3E6F: data = 12'h502;
        15'h3E70: data = 12'h510;
        15'h3E71: data = 12'h524;
        15'h3E72: data = 12'h539;
        15'h3E73: data = 12'h549;
        15'h3E74: data = 12'h55C;
        15'h3E75: data = 12'h56A;
        15'h3E76: data = 12'h581;
        15'h3E77: data = 12'h593;
        15'h3E78: data = 12'h5A7;
        15'h3E79: data = 12'h5BA;
        15'h3E7A: data = 12'h5C8;
        15'h3E7B: data = 12'h5DA;
        15'h3E7C: data = 12'h5F1;
        15'h3E7D: data = 12'h600;
        15'h3E7E: data = 12'h60C;
        15'h3E7F: data = 12'h621;
        15'h3E80: data = 12'h634;
        15'h3E81: data = 12'h645;
        15'h3E82: data = 12'h657;
        15'h3E83: data = 12'h66B;
        15'h3E84: data = 12'h67A;
        15'h3E85: data = 12'h686;
        15'h3E86: data = 12'h699;
        15'h3E87: data = 12'h6A7;
        15'h3E88: data = 12'h6BA;
        15'h3E89: data = 12'h6C5;
        15'h3E8A: data = 12'h6D5;
        15'h3E8B: data = 12'h6DF;
        15'h3E8C: data = 12'h6F0;
        15'h3E8D: data = 12'h6FD;
        15'h3E8E: data = 12'h70D;
        15'h3E8F: data = 12'h714;
        15'h3E90: data = 12'h724;
        15'h3E91: data = 12'h735;
        15'h3E92: data = 12'h73A;
        15'h3E93: data = 12'h747;
        15'h3E94: data = 12'h74E;
        15'h3E95: data = 12'h75D;
        15'h3E96: data = 12'h765;
        15'h3E97: data = 12'h775;
        15'h3E98: data = 12'h77A;
        15'h3E99: data = 12'h78E;
        15'h3E9A: data = 12'h793;
        15'h3E9B: data = 12'h79B;
        15'h3E9C: data = 12'h7A2;
        15'h3E9D: data = 12'h7B1;
        15'h3E9E: data = 12'h7B5;
        15'h3E9F: data = 12'h7B9;
        15'h3EA0: data = 12'h7C3;
        15'h3EA1: data = 12'h7CA;
        15'h3EA2: data = 12'h7D0;
        15'h3EA3: data = 12'h7D7;
        15'h3EA4: data = 12'h7E5;
        15'h3EA5: data = 12'h7E6;
        15'h3EA6: data = 12'h7EE;
        15'h3EA7: data = 12'h7EF;
        15'h3EA8: data = 12'h7FB;
        15'h3EA9: data = 12'h7FC;
        15'h3EAA: data = 12'h7FC;
        15'h3EAB: data = 12'h804;
        15'h3EAC: data = 12'h6CA;
        15'h3EAD: data = 12'h085;
        15'h3EAE: data = 12'h092;
        15'h3EAF: data = 12'h093;
        15'h3EB0: data = 12'h093;
        15'h3EB1: data = 12'h09C;
        15'h3EB2: data = 12'h09F;
        15'h3EB3: data = 12'h0AA;
        15'h3EB4: data = 12'h0AB;
        15'h3EB5: data = 12'h0AC;
        15'h3EB6: data = 12'h0B4;
        15'h3EB7: data = 12'h0B9;
        15'h3EB8: data = 12'h0BB;
        15'h3EB9: data = 12'h0C1;
        15'h3EBA: data = 12'h0CB;
        15'h3EBB: data = 12'h0CD;
        15'h3EBC: data = 12'h0D1;
        15'h3EBD: data = 12'h0D6;
        15'h3EBE: data = 12'h0D8;
        15'h3EBF: data = 12'h0D6;
        15'h3EC0: data = 12'h0D5;
        15'h3EC1: data = 12'h0CE;
        15'h3EC2: data = 12'h0CA;
        15'h3EC3: data = 12'h0C8;
        15'h3EC4: data = 12'h0C4;
        15'h3EC5: data = 12'h0BC;
        15'h3EC6: data = 12'h0B9;
        15'h3EC7: data = 12'h0B3;
        15'h3EC8: data = 12'h0AF;
        15'h3EC9: data = 12'h0B0;
        15'h3ECA: data = 12'h0A9;
        15'h3ECB: data = 12'h0B2;
        15'h3ECC: data = 12'h0B0;
        15'h3ECD: data = 12'h0B5;
        15'h3ECE: data = 12'h0AD;
        15'h3ECF: data = 12'h0A5;
        15'h3ED0: data = 12'h0A5;
        15'h3ED1: data = 12'h09C;
        15'h3ED2: data = 12'h08A;
        15'h3ED3: data = 12'h07C;
        15'h3ED4: data = 12'h072;
        15'h3ED5: data = 12'h074;
        15'h3ED6: data = 12'h06F;
        15'h3ED7: data = 12'h06D;
        15'h3ED8: data = 12'h06B;
        15'h3ED9: data = 12'h069;
        15'h3EDA: data = 12'h060;
        15'h3EDB: data = 12'h054;
        15'h3EDC: data = 12'h042;
        15'h3EDD: data = 12'h7BB;
        15'h3EDE: data = 12'h7B1;
        15'h3EDF: data = 12'h7A6;
        15'h3EE0: data = 12'h7A7;
        15'h3EE1: data = 12'h79B;
        15'h3EE2: data = 12'h794;
        15'h3EE3: data = 12'h787;
        15'h3EE4: data = 12'h77B;
        15'h3EE5: data = 12'h769;
        15'h3EE6: data = 12'h758;
        15'h3EE7: data = 12'h741;
        15'h3EE8: data = 12'h736;
        15'h3EE9: data = 12'h72E;
        15'h3EEA: data = 12'h726;
        15'h3EEB: data = 12'h71B;
        15'h3EEC: data = 12'h712;
        15'h3EED: data = 12'h70B;
        15'h3EEE: data = 12'h6FC;
        15'h3EEF: data = 12'h6E8;
        15'h3EF0: data = 12'h6DB;
        15'h3EF1: data = 12'h6C5;
        15'h3EF2: data = 12'h6B4;
        15'h3EF3: data = 12'h6A2;
        15'h3EF4: data = 12'h695;
        15'h3EF5: data = 12'h689;
        15'h3EF6: data = 12'h67B;
        15'h3EF7: data = 12'h672;
        15'h3EF8: data = 12'h668;
        15'h3EF9: data = 12'h657;
        15'h3EFA: data = 12'h645;
        15'h3EFB: data = 12'h632;
        15'h3EFC: data = 12'h62A;
        15'h3EFD: data = 12'h610;
        15'h3EFE: data = 12'h5F9;
        15'h3EFF: data = 12'h5E8;
        15'h3F00: data = 12'h5D0;
        15'h3F01: data = 12'h5C0;
        15'h3F02: data = 12'h5B3;
        15'h3F03: data = 12'h59F;
        15'h3F04: data = 12'h591;
        15'h3F05: data = 12'h582;
        15'h3F06: data = 12'h574;
        15'h3F07: data = 12'h564;
        15'h3F08: data = 12'h552;
        15'h3F09: data = 12'h542;
        15'h3F0A: data = 12'h52D;
        15'h3F0B: data = 12'h516;
        15'h3F0C: data = 12'h508;
        15'h3F0D: data = 12'h4F4;
        15'h3F0E: data = 12'h4DA;
        15'h3F0F: data = 12'h4C2;
        15'h3F10: data = 12'h4B1;
        15'h3F11: data = 12'h495;
        15'h3F12: data = 12'h47D;
        15'h3F13: data = 12'h469;
        15'h3F14: data = 12'h44F;
        15'h3F15: data = 12'h440;
        15'h3F16: data = 12'h429;
        15'h3F17: data = 12'h413;
        15'h3F18: data = 12'h3FD;
        15'h3F19: data = 12'h3E9;
        15'h3F1A: data = 12'h3CE;
        15'h3F1B: data = 12'h3BC;
        15'h3F1C: data = 12'h3A9;
        15'h3F1D: data = 12'h392;
        15'h3F1E: data = 12'h37F;
        15'h3F1F: data = 12'h36C;
        15'h3F20: data = 12'h355;
        15'h3F21: data = 12'h33F;
        15'h3F22: data = 12'h32A;
        15'h3F23: data = 12'h315;
        15'h3F24: data = 12'h2FC;
        15'h3F25: data = 12'h2E8;
        15'h3F26: data = 12'h2D6;
        15'h3F27: data = 12'h2BF;
        15'h3F28: data = 12'h2A8;
        15'h3F29: data = 12'h28F;
        15'h3F2A: data = 12'h27E;
        15'h3F2B: data = 12'h267;
        15'h3F2C: data = 12'h24A;
        15'h3F2D: data = 12'h236;
        15'h3F2E: data = 12'h21E;
        15'h3F2F: data = 12'h205;
        15'h3F30: data = 12'h1F1;
        15'h3F31: data = 12'h1DA;
        15'h3F32: data = 12'h1C4;
        15'h3F33: data = 12'h1AA;
        15'h3F34: data = 12'h193;
        15'h3F35: data = 12'h17D;
        15'h3F36: data = 12'h165;
        15'h3F37: data = 12'h151;
        15'h3F38: data = 12'h139;
        15'h3F39: data = 12'h11F;
        15'h3F3A: data = 12'h109;
        15'h3F3B: data = 12'h0F4;
        15'h3F3C: data = 12'h0DA;
        15'h3F3D: data = 12'h0BF;
        15'h3F3E: data = 12'h0A9;
        15'h3F3F: data = 12'h090;
        15'h3F40: data = 12'h07E;
        15'h3F41: data = 12'h065;
        15'h3F42: data = 12'h04D;
        15'h3F43: data = 12'h7E0;
        15'h3F44: data = 12'h7CD;
        15'h3F45: data = 12'h7B8;
        15'h3F46: data = 12'h7A3;
        15'h3F47: data = 12'h78E;
        15'h3F48: data = 12'h775;
        15'h3F49: data = 12'h75A;
        15'h3F4A: data = 12'h747;
        15'h3F4B: data = 12'h734;
        15'h3F4C: data = 12'h71A;
        15'h3F4D: data = 12'h703;
        15'h3F4E: data = 12'h6E8;
        15'h3F4F: data = 12'h6DB;
        15'h3F50: data = 12'h6C3;
        15'h3F51: data = 12'h6AF;
        15'h3F52: data = 12'h690;
        15'h3F53: data = 12'h67F;
        15'h3F54: data = 12'h665;
        15'h3F55: data = 12'h650;
        15'h3F56: data = 12'h63B;
        15'h3F57: data = 12'h625;
        15'h3F58: data = 12'h611;
        15'h3F59: data = 12'h5F6;
        15'h3F5A: data = 12'h5E1;
        15'h3F5B: data = 12'h5CA;
        15'h3F5C: data = 12'h5B4;
        15'h3F5D: data = 12'h597;
        15'h3F5E: data = 12'h580;
        15'h3F5F: data = 12'h56C;
        15'h3F60: data = 12'h55A;
        15'h3F61: data = 12'h547;
        15'h3F62: data = 12'h531;
        15'h3F63: data = 12'h519;
        15'h3F64: data = 12'h505;
        15'h3F65: data = 12'h4F1;
        15'h3F66: data = 12'h4DE;
        15'h3F67: data = 12'h4C7;
        15'h3F68: data = 12'h4B5;
        15'h3F69: data = 12'h49F;
        15'h3F6A: data = 12'h490;
        15'h3F6B: data = 12'h47B;
        15'h3F6C: data = 12'h46A;
        15'h3F6D: data = 12'h45A;
        15'h3F6E: data = 12'h44B;
        15'h3F6F: data = 12'h43A;
        15'h3F70: data = 12'h42A;
        15'h3F71: data = 12'h416;
        15'h3F72: data = 12'h407;
        15'h3F73: data = 12'h3F8;
        15'h3F74: data = 12'h3EA;
        15'h3F75: data = 12'h3D0;
        15'h3F76: data = 12'h3C5;
        15'h3F77: data = 12'h3AD;
        15'h3F78: data = 12'h399;
        15'h3F79: data = 12'h38E;
        15'h3F7A: data = 12'h377;
        15'h3F7B: data = 12'h366;
        15'h3F7C: data = 12'h352;
        15'h3F7D: data = 12'h33F;
        15'h3F7E: data = 12'h32D;
        15'h3F7F: data = 12'h31C;
        15'h3F80: data = 12'h30F;
        15'h3F81: data = 12'h2FF;
        15'h3F82: data = 12'h2F0;
        15'h3F83: data = 12'h2DD;
        15'h3F84: data = 12'h2D6;
        15'h3F85: data = 12'h2D1;
        15'h3F86: data = 12'h2C7;
        15'h3F87: data = 12'h2BB;
        15'h3F88: data = 12'h2AB;
        15'h3F89: data = 12'h29C;
        15'h3F8A: data = 12'h293;
        15'h3F8B: data = 12'h287;
        15'h3F8C: data = 12'h27B;
        15'h3F8D: data = 12'h269;
        15'h3F8E: data = 12'h25D;
        15'h3F8F: data = 12'h24C;
        15'h3F90: data = 12'h23D;
        15'h3F91: data = 12'h22F;
        15'h3F92: data = 12'h221;
        15'h3F93: data = 12'h218;
        15'h3F94: data = 12'h211;
        15'h3F95: data = 12'h20E;
        15'h3F96: data = 12'h203;
        15'h3F97: data = 12'h1FB;
        15'h3F98: data = 12'h1F6;
        15'h3F99: data = 12'h1F1;
        15'h3F9A: data = 12'h1ED;
        15'h3F9B: data = 12'h1DE;
        15'h3F9C: data = 12'h1D4;
        15'h3F9D: data = 12'h1CA;
        15'h3F9E: data = 12'h1C2;
        15'h3F9F: data = 12'h1BD;
        15'h3FA0: data = 12'h1B4;
        15'h3FA1: data = 12'h1A6;
        15'h3FA2: data = 12'h198;
        15'h3FA3: data = 12'h193;
        15'h3FA4: data = 12'h192;
        15'h3FA5: data = 12'h18E;
        15'h3FA6: data = 12'h18D;
        15'h3FA7: data = 12'h186;
        15'h3FA8: data = 12'h18B;
        15'h3FA9: data = 12'h186;
        15'h3FAA: data = 12'h186;
        15'h3FAB: data = 12'h17E;
        15'h3FAC: data = 12'h17E;
        15'h3FAD: data = 12'h175;
        15'h3FAE: data = 12'h171;
        15'h3FAF: data = 12'h16D;
        15'h3FB0: data = 12'h165;
        15'h3FB1: data = 12'h15F;
        15'h3FB2: data = 12'h15D;
        15'h3FB3: data = 12'h15D;
        15'h3FB4: data = 12'h158;
        15'h3FB5: data = 12'h159;
        15'h3FB6: data = 12'h15C;
        15'h3FB7: data = 12'h161;
        15'h3FB8: data = 12'h166;
        15'h3FB9: data = 12'h166;
        15'h3FBA: data = 12'h169;
        15'h3FBB: data = 12'h171;
        15'h3FBC: data = 12'h16E;
        15'h3FBD: data = 12'h16C;
        15'h3FBE: data = 12'h16A;
        15'h3FBF: data = 12'h168;
        15'h3FC0: data = 12'h169;
        15'h3FC1: data = 12'h166;
        15'h3FC2: data = 12'h16C;
        15'h3FC3: data = 12'h16C;
        15'h3FC4: data = 12'h16D;
        15'h3FC5: data = 12'h177;
        15'h3FC6: data = 12'h181;
        15'h3FC7: data = 12'h185;
        15'h3FC8: data = 12'h190;
        15'h3FC9: data = 12'h197;
        15'h3FCA: data = 12'h199;
        15'h3FCB: data = 12'h1A7;
        15'h3FCC: data = 12'h1AC;
        15'h3FCD: data = 12'h1B0;
        15'h3FCE: data = 12'h1B3;
        15'h3FCF: data = 12'h1B6;
        15'h3FD0: data = 12'h1B6;
        15'h3FD1: data = 12'h1BB;
        15'h3FD2: data = 12'h1C0;
        15'h3FD3: data = 12'h1C7;
        15'h3FD4: data = 12'h1D2;
        15'h3FD5: data = 12'h1DB;
        15'h3FD6: data = 12'h1E8;
        15'h3FD7: data = 12'h1F4;
        15'h3FD8: data = 12'h1FF;
        15'h3FD9: data = 12'h20B;
        15'h3FDA: data = 12'h21D;
        15'h3FDB: data = 12'h21F;
        15'h3FDC: data = 12'h22F;
        15'h3FDD: data = 12'h23A;
        15'h3FDE: data = 12'h248;
        15'h3FDF: data = 12'h24C;
        15'h3FE0: data = 12'h25B;
        15'h3FE1: data = 12'h263;
        15'h3FE2: data = 12'h26D;
        15'h3FE3: data = 12'h270;
        15'h3FE4: data = 12'h27E;
        15'h3FE5: data = 12'h28B;
        15'h3FE6: data = 12'h290;
        15'h3FE7: data = 12'h2A3;
        15'h3FE8: data = 12'h2AE;
        15'h3FE9: data = 12'h2C3;
        15'h3FEA: data = 12'h2D5;
        15'h3FEB: data = 12'h2DE;
        15'h3FEC: data = 12'h2F2;
        15'h3FED: data = 12'h306;
        15'h3FEE: data = 12'h31A;
        15'h3FEF: data = 12'h32A;
        15'h3FF0: data = 12'h339;
        15'h3FF1: data = 12'h344;
        15'h3FF2: data = 12'h356;
        15'h3FF3: data = 12'h365;
        15'h3FF4: data = 12'h371;
        15'h3FF5: data = 12'h37E;
        15'h3FF6: data = 12'h38E;
        15'h3FF7: data = 12'h396;
        15'h3FF8: data = 12'h3AA;
        15'h3FF9: data = 12'h3B6;
        15'h3FFA: data = 12'h3C4;
        15'h3FFB: data = 12'h3DE;
        15'h3FFC: data = 12'h3EC;
        15'h3FFD: data = 12'h400;
        15'h3FFE: data = 12'h417;
        15'h3FFF: data = 12'h42B;
        15'h4000: data = 12'h444;
        15'h4001: data = 12'h455;
        15'h4002: data = 12'h469;
        15'h4003: data = 12'h480;
        15'h4004: data = 12'h494;
        15'h4005: data = 12'h4AC;
        15'h4006: data = 12'h4B8;
        15'h4007: data = 12'h4D0;
        15'h4008: data = 12'h4E8;
        15'h4009: data = 12'h4FA;
        15'h400A: data = 12'h50C;
        15'h400B: data = 12'h519;
        15'h400C: data = 12'h526;
        15'h400D: data = 12'h53B;
        15'h400E: data = 12'h552;
        15'h400F: data = 12'h563;
        15'h4010: data = 12'h577;
        15'h4011: data = 12'h58A;
        15'h4012: data = 12'h5A1;
        15'h4013: data = 12'h5B8;
        15'h4014: data = 12'h5CE;
        15'h4015: data = 12'h5E7;
        15'h4016: data = 12'h601;
        15'h4017: data = 12'h619;
        15'h4018: data = 12'h635;
        15'h4019: data = 12'h64A;
        15'h401A: data = 12'h660;
        15'h401B: data = 12'h677;
        15'h401C: data = 12'h692;
        15'h401D: data = 12'h6A1;
        15'h401E: data = 12'h6B5;
        15'h401F: data = 12'h6CF;
        15'h4020: data = 12'h6E0;
        15'h4021: data = 12'h6F6;
        15'h4022: data = 12'h708;
        15'h4023: data = 12'h71C;
        15'h4024: data = 12'h739;
        15'h4025: data = 12'h744;
        15'h4026: data = 12'h75A;
        15'h4027: data = 12'h776;
        15'h4028: data = 12'h790;
        15'h4029: data = 12'h7A3;
        15'h402A: data = 12'h7BD;
        15'h402B: data = 12'h7D6;
        15'h402C: data = 12'h7EA;
        15'h402D: data = 12'h804;
        15'h402E: data = 12'h076;
        15'h402F: data = 12'h08C;
        15'h4030: data = 12'h0A1;
        15'h4031: data = 12'h0B8;
        15'h4032: data = 12'h0D3;
        15'h4033: data = 12'h0E8;
        15'h4034: data = 12'h101;
        15'h4035: data = 12'h113;
        15'h4036: data = 12'h128;
        15'h4037: data = 12'h145;
        15'h4038: data = 12'h157;
        15'h4039: data = 12'h16D;
        15'h403A: data = 12'h182;
        15'h403B: data = 12'h199;
        15'h403C: data = 12'h1AF;
        15'h403D: data = 12'h1BD;
        15'h403E: data = 12'h1D7;
        15'h403F: data = 12'h1ED;
        15'h4040: data = 12'h205;
        15'h4041: data = 12'h218;
        15'h4042: data = 12'h232;
        15'h4043: data = 12'h246;
        15'h4044: data = 12'h25F;
        15'h4045: data = 12'h276;
        15'h4046: data = 12'h290;
        15'h4047: data = 12'h2A8;
        15'h4048: data = 12'h2C2;
        15'h4049: data = 12'h2DC;
        15'h404A: data = 12'h2F2;
        15'h404B: data = 12'h30C;
        15'h404C: data = 12'h327;
        15'h404D: data = 12'h33C;
        15'h404E: data = 12'h34F;
        15'h404F: data = 12'h36C;
        15'h4050: data = 12'h381;
        15'h4051: data = 12'h39A;
        15'h4052: data = 12'h3AD;
        15'h4053: data = 12'h3C3;
        15'h4054: data = 12'h3D6;
        15'h4055: data = 12'h3F4;
        15'h4056: data = 12'h405;
        15'h4057: data = 12'h416;
        15'h4058: data = 12'h42E;
        15'h4059: data = 12'h443;
        15'h405A: data = 12'h452;
        15'h405B: data = 12'h467;
        15'h405C: data = 12'h47C;
        15'h405D: data = 12'h493;
        15'h405E: data = 12'h4A6;
        15'h405F: data = 12'h4B5;
        15'h4060: data = 12'h4C5;
        15'h4061: data = 12'h4DA;
        15'h4062: data = 12'h4ED;
        15'h4063: data = 12'h505;
        15'h4064: data = 12'h511;
        15'h4065: data = 12'h528;
        15'h4066: data = 12'h53B;
        15'h4067: data = 12'h54B;
        15'h4068: data = 12'h555;
        15'h4069: data = 12'h569;
        15'h406A: data = 12'h57E;
        15'h406B: data = 12'h58F;
        15'h406C: data = 12'h5A4;
        15'h406D: data = 12'h5B5;
        15'h406E: data = 12'h5C5;
        15'h406F: data = 12'h5D9;
        15'h4070: data = 12'h5ED;
        15'h4071: data = 12'h5FD;
        15'h4072: data = 12'h60F;
        15'h4073: data = 12'h61E;
        15'h4074: data = 12'h632;
        15'h4075: data = 12'h642;
        15'h4076: data = 12'h656;
        15'h4077: data = 12'h666;
        15'h4078: data = 12'h674;
        15'h4079: data = 12'h688;
        15'h407A: data = 12'h699;
        15'h407B: data = 12'h6A8;
        15'h407C: data = 12'h6B8;
        15'h407D: data = 12'h6C3;
        15'h407E: data = 12'h6D6;
        15'h407F: data = 12'h6E0;
        15'h4080: data = 12'h6EE;
        15'h4081: data = 12'h6FF;
        15'h4082: data = 12'h70D;
        15'h4083: data = 12'h717;
        15'h4084: data = 12'h725;
        15'h4085: data = 12'h735;
        15'h4086: data = 12'h73D;
        15'h4087: data = 12'h748;
        15'h4088: data = 12'h750;
        15'h4089: data = 12'h75F;
        15'h408A: data = 12'h766;
        15'h408B: data = 12'h776;
        15'h408C: data = 12'h77F;
        15'h408D: data = 12'h78E;
        15'h408E: data = 12'h797;
        15'h408F: data = 12'h79A;
        15'h4090: data = 12'h7A0;
        15'h4091: data = 12'h7AD;
        15'h4092: data = 12'h7B4;
        15'h4093: data = 12'h7C0;
        15'h4094: data = 12'h7C4;
        15'h4095: data = 12'h7CC;
        15'h4096: data = 12'h7D3;
        15'h4097: data = 12'h7D9;
        15'h4098: data = 12'h7E5;
        15'h4099: data = 12'h7EA;
        15'h409A: data = 12'h7EF;
        15'h409B: data = 12'h7F4;
        15'h409C: data = 12'h7F9;
        15'h409D: data = 12'h800;
        15'h409E: data = 12'h7FE;
        15'h409F: data = 12'h806;
        15'h40A0: data = 12'h73E;
        15'h40A1: data = 12'h082;
        15'h40A2: data = 12'h08F;
        15'h40A3: data = 12'h096;
        15'h40A4: data = 12'h096;
        15'h40A5: data = 12'h09F;
        15'h40A6: data = 12'h0A0;
        15'h40A7: data = 12'h0A8;
        15'h40A8: data = 12'h0AB;
        15'h40A9: data = 12'h0AB;
        15'h40AA: data = 12'h0B6;
        15'h40AB: data = 12'h0B4;
        15'h40AC: data = 12'h0B9;
        15'h40AD: data = 12'h0BE;
        15'h40AE: data = 12'h0C9;
        15'h40AF: data = 12'h0CB;
        15'h40B0: data = 12'h0CF;
        15'h40B1: data = 12'h0D4;
        15'h40B2: data = 12'h0D2;
        15'h40B3: data = 12'h0D5;
        15'h40B4: data = 12'h0D5;
        15'h40B5: data = 12'h0CD;
        15'h40B6: data = 12'h0CE;
        15'h40B7: data = 12'h0CA;
        15'h40B8: data = 12'h0C7;
        15'h40B9: data = 12'h0C1;
        15'h40BA: data = 12'h0B7;
        15'h40BB: data = 12'h0B2;
        15'h40BC: data = 12'h0AA;
        15'h40BD: data = 12'h0AF;
        15'h40BE: data = 12'h0A8;
        15'h40BF: data = 12'h0AB;
        15'h40C0: data = 12'h0AF;
        15'h40C1: data = 12'h0B5;
        15'h40C2: data = 12'h0AD;
        15'h40C3: data = 12'h0A6;
        15'h40C4: data = 12'h0A4;
        15'h40C5: data = 12'h099;
        15'h40C6: data = 12'h08E;
        15'h40C7: data = 12'h07E;
        15'h40C8: data = 12'h072;
        15'h40C9: data = 12'h076;
        15'h40CA: data = 12'h06C;
        15'h40CB: data = 12'h06C;
        15'h40CC: data = 12'h06C;
        15'h40CD: data = 12'h06A;
        15'h40CE: data = 12'h062;
        15'h40CF: data = 12'h054;
        15'h40D0: data = 12'h044;
        15'h40D1: data = 12'h7BE;
        15'h40D2: data = 12'h7B2;
        15'h40D3: data = 12'h7A6;
        15'h40D4: data = 12'h7A1;
        15'h40D5: data = 12'h797;
        15'h40D6: data = 12'h792;
        15'h40D7: data = 12'h78B;
        15'h40D8: data = 12'h77B;
        15'h40D9: data = 12'h768;
        15'h40DA: data = 12'h759;
        15'h40DB: data = 12'h740;
        15'h40DC: data = 12'h736;
        15'h40DD: data = 12'h72E;
        15'h40DE: data = 12'h727;
        15'h40DF: data = 12'h71A;
        15'h40E0: data = 12'h712;
        15'h40E1: data = 12'h70A;
        15'h40E2: data = 12'h6FA;
        15'h40E3: data = 12'h6EA;
        15'h40E4: data = 12'h6DA;
        15'h40E5: data = 12'h6C6;
        15'h40E6: data = 12'h6B3;
        15'h40E7: data = 12'h6A4;
        15'h40E8: data = 12'h695;
        15'h40E9: data = 12'h688;
        15'h40EA: data = 12'h67F;
        15'h40EB: data = 12'h673;
        15'h40EC: data = 12'h666;
        15'h40ED: data = 12'h657;
        15'h40EE: data = 12'h646;
        15'h40EF: data = 12'h633;
        15'h40F0: data = 12'h62A;
        15'h40F1: data = 12'h611;
        15'h40F2: data = 12'h5FE;
        15'h40F3: data = 12'h5E7;
        15'h40F4: data = 12'h5CD;
        15'h40F5: data = 12'h5BC;
        15'h40F6: data = 12'h5AF;
        15'h40F7: data = 12'h5A0;
        15'h40F8: data = 12'h58F;
        15'h40F9: data = 12'h580;
        15'h40FA: data = 12'h56F;
        15'h40FB: data = 12'h564;
        15'h40FC: data = 12'h555;
        15'h40FD: data = 12'h542;
        15'h40FE: data = 12'h52D;
        15'h40FF: data = 12'h518;
        15'h4100: data = 12'h507;
        15'h4101: data = 12'h4F3;
        15'h4102: data = 12'h4DB;
        15'h4103: data = 12'h4C7;
        15'h4104: data = 12'h4B2;
        15'h4105: data = 12'h497;
        15'h4106: data = 12'h47D;
        15'h4107: data = 12'h466;
        15'h4108: data = 12'h44F;
        15'h4109: data = 12'h43E;
        15'h410A: data = 12'h429;
        15'h410B: data = 12'h413;
        15'h410C: data = 12'h3FE;
        15'h410D: data = 12'h3E8;
        15'h410E: data = 12'h3D0;
        15'h410F: data = 12'h3C0;
        15'h4110: data = 12'h3A9;
        15'h4111: data = 12'h38E;
        15'h4112: data = 12'h381;
        15'h4113: data = 12'h36A;
        15'h4114: data = 12'h358;
        15'h4115: data = 12'h342;
        15'h4116: data = 12'h32B;
        15'h4117: data = 12'h318;
        15'h4118: data = 12'h2FE;
        15'h4119: data = 12'h2EA;
        15'h411A: data = 12'h2D9;
        15'h411B: data = 12'h2C3;
        15'h411C: data = 12'h2A5;
        15'h411D: data = 12'h292;
        15'h411E: data = 12'h280;
        15'h411F: data = 12'h264;
        15'h4120: data = 12'h24A;
        15'h4121: data = 12'h236;
        15'h4122: data = 12'h21C;
        15'h4123: data = 12'h206;
        15'h4124: data = 12'h1F0;
        15'h4125: data = 12'h1D8;
        15'h4126: data = 12'h1C4;
        15'h4127: data = 12'h1AC;
        15'h4128: data = 12'h192;
        15'h4129: data = 12'h17B;
        15'h412A: data = 12'h168;
        15'h412B: data = 12'h150;
        15'h412C: data = 12'h137;
        15'h412D: data = 12'h11C;
        15'h412E: data = 12'h108;
        15'h412F: data = 12'h0F5;
        15'h4130: data = 12'h0D8;
        15'h4131: data = 12'h0C2;
        15'h4132: data = 12'h0A8;
        15'h4133: data = 12'h091;
        15'h4134: data = 12'h07B;
        15'h4135: data = 12'h062;
        15'h4136: data = 12'h04C;
        15'h4137: data = 12'h7E3;
        15'h4138: data = 12'h7CC;
        15'h4139: data = 12'h7B6;
        15'h413A: data = 12'h7A3;
        15'h413B: data = 12'h78E;
        15'h413C: data = 12'h777;
        15'h413D: data = 12'h759;
        15'h413E: data = 12'h748;
        15'h413F: data = 12'h736;
        15'h4140: data = 12'h71F;
        15'h4141: data = 12'h705;
        15'h4142: data = 12'h6E8;
        15'h4143: data = 12'h6DA;
        15'h4144: data = 12'h6C2;
        15'h4145: data = 12'h6AA;
        15'h4146: data = 12'h68F;
        15'h4147: data = 12'h67E;
        15'h4148: data = 12'h665;
        15'h4149: data = 12'h651;
        15'h414A: data = 12'h63B;
        15'h414B: data = 12'h626;
        15'h414C: data = 12'h60E;
        15'h414D: data = 12'h5F0;
        15'h414E: data = 12'h5E0;
        15'h414F: data = 12'h5CA;
        15'h4150: data = 12'h5B3;
        15'h4151: data = 12'h59B;
        15'h4152: data = 12'h582;
        15'h4153: data = 12'h56D;
        15'h4154: data = 12'h55C;
        15'h4155: data = 12'h544;
        15'h4156: data = 12'h52C;
        15'h4157: data = 12'h51A;
        15'h4158: data = 12'h504;
        15'h4159: data = 12'h4F3;
        15'h415A: data = 12'h4DA;
        15'h415B: data = 12'h4CC;
        15'h415C: data = 12'h4B6;
        15'h415D: data = 12'h4A2;
        15'h415E: data = 12'h492;
        15'h415F: data = 12'h47F;
        15'h4160: data = 12'h46C;
        15'h4161: data = 12'h45D;
        15'h4162: data = 12'h44B;
        15'h4163: data = 12'h43C;
        15'h4164: data = 12'h42C;
        15'h4165: data = 12'h419;
        15'h4166: data = 12'h409;
        15'h4167: data = 12'h3F8;
        15'h4168: data = 12'h3E9;
        15'h4169: data = 12'h3D3;
        15'h416A: data = 12'h3C2;
        15'h416B: data = 12'h3AC;
        15'h416C: data = 12'h39B;
        15'h416D: data = 12'h38C;
        15'h416E: data = 12'h373;
        15'h416F: data = 12'h363;
        15'h4170: data = 12'h34E;
        15'h4171: data = 12'h341;
        15'h4172: data = 12'h32C;
        15'h4173: data = 12'h31D;
        15'h4174: data = 12'h30E;
        15'h4175: data = 12'h2FF;
        15'h4176: data = 12'h2F4;
        15'h4177: data = 12'h2E4;
        15'h4178: data = 12'h2D9;
        15'h4179: data = 12'h2D4;
        15'h417A: data = 12'h2C8;
        15'h417B: data = 12'h2BE;
        15'h417C: data = 12'h2AD;
        15'h417D: data = 12'h29F;
        15'h417E: data = 12'h295;
        15'h417F: data = 12'h285;
        15'h4180: data = 12'h27C;
        15'h4181: data = 12'h268;
        15'h4182: data = 12'h258;
        15'h4183: data = 12'h248;
        15'h4184: data = 12'h239;
        15'h4185: data = 12'h22B;
        15'h4186: data = 12'h21F;
        15'h4187: data = 12'h215;
        15'h4188: data = 12'h211;
        15'h4189: data = 12'h20C;
        15'h418A: data = 12'h206;
        15'h418B: data = 12'h1FC;
        15'h418C: data = 12'h1F8;
        15'h418D: data = 12'h1EF;
        15'h418E: data = 12'h1E8;
        15'h418F: data = 12'h1DE;
        15'h4190: data = 12'h1D0;
        15'h4191: data = 12'h1C8;
        15'h4192: data = 12'h1C0;
        15'h4193: data = 12'h1B6;
        15'h4194: data = 12'h1AB;
        15'h4195: data = 12'h1A3;
        15'h4196: data = 12'h19B;
        15'h4197: data = 12'h191;
        15'h4198: data = 12'h18F;
        15'h4199: data = 12'h18F;
        15'h419A: data = 12'h18C;
        15'h419B: data = 12'h18A;
        15'h419C: data = 12'h18B;
        15'h419D: data = 12'h189;
        15'h419E: data = 12'h187;
        15'h419F: data = 12'h17D;
        15'h41A0: data = 12'h17E;
        15'h41A1: data = 12'h172;
        15'h41A2: data = 12'h16C;
        15'h41A3: data = 12'h16B;
        15'h41A4: data = 12'h160;
        15'h41A5: data = 12'h15E;
        15'h41A6: data = 12'h15B;
        15'h41A7: data = 12'h15E;
        15'h41A8: data = 12'h157;
        15'h41A9: data = 12'h15A;
        15'h41AA: data = 12'h15E;
        15'h41AB: data = 12'h164;
        15'h41AC: data = 12'h168;
        15'h41AD: data = 12'h169;
        15'h41AE: data = 12'h16B;
        15'h41AF: data = 12'h16F;
        15'h41B0: data = 12'h170;
        15'h41B1: data = 12'h16B;
        15'h41B2: data = 12'h167;
        15'h41B3: data = 12'h165;
        15'h41B4: data = 12'h168;
        15'h41B5: data = 12'h164;
        15'h41B6: data = 12'h16D;
        15'h41B7: data = 12'h16C;
        15'h41B8: data = 12'h172;
        15'h41B9: data = 12'h174;
        15'h41BA: data = 12'h185;
        15'h41BB: data = 12'h189;
        15'h41BC: data = 12'h191;
        15'h41BD: data = 12'h197;
        15'h41BE: data = 12'h19E;
        15'h41BF: data = 12'h1A9;
        15'h41C0: data = 12'h1AC;
        15'h41C1: data = 12'h1B0;
        15'h41C2: data = 12'h1B5;
        15'h41C3: data = 12'h1B6;
        15'h41C4: data = 12'h1B9;
        15'h41C5: data = 12'h1BF;
        15'h41C6: data = 12'h1C4;
        15'h41C7: data = 12'h1C9;
        15'h41C8: data = 12'h1CF;
        15'h41C9: data = 12'h1D7;
        15'h41CA: data = 12'h1E8;
        15'h41CB: data = 12'h1F7;
        15'h41CC: data = 12'h200;
        15'h41CD: data = 12'h20D;
        15'h41CE: data = 12'h21F;
        15'h41CF: data = 12'h222;
        15'h41D0: data = 12'h233;
        15'h41D1: data = 12'h23B;
        15'h41D2: data = 12'h249;
        15'h41D3: data = 12'h24D;
        15'h41D4: data = 12'h258;
        15'h41D5: data = 12'h263;
        15'h41D6: data = 12'h26D;
        15'h41D7: data = 12'h270;
        15'h41D8: data = 12'h27A;
        15'h41D9: data = 12'h289;
        15'h41DA: data = 12'h28F;
        15'h41DB: data = 12'h2A1;
        15'h41DC: data = 12'h2AF;
        15'h41DD: data = 12'h2C5;
        15'h41DE: data = 12'h2D9;
        15'h41DF: data = 12'h2DF;
        15'h41E0: data = 12'h2F6;
        15'h41E1: data = 12'h307;
        15'h41E2: data = 12'h318;
        15'h41E3: data = 12'h327;
        15'h41E4: data = 12'h338;
        15'h41E5: data = 12'h344;
        15'h41E6: data = 12'h355;
        15'h41E7: data = 12'h361;
        15'h41E8: data = 12'h370;
        15'h41E9: data = 12'h37A;
        15'h41EA: data = 12'h38F;
        15'h41EB: data = 12'h396;
        15'h41EC: data = 12'h3A9;
        15'h41ED: data = 12'h3B7;
        15'h41EE: data = 12'h3C6;
        15'h41EF: data = 12'h3DE;
        15'h41F0: data = 12'h3ED;
        15'h41F1: data = 12'h3FE;
        15'h41F2: data = 12'h41B;
        15'h41F3: data = 12'h42E;
        15'h41F4: data = 12'h444;
        15'h41F5: data = 12'h45C;
        15'h41F6: data = 12'h46D;
        15'h41F7: data = 12'h484;
        15'h41F8: data = 12'h495;
        15'h41F9: data = 12'h4AA;
        15'h41FA: data = 12'h4BC;
        15'h41FB: data = 12'h4D0;
        15'h41FC: data = 12'h4E5;
        15'h41FD: data = 12'h4F8;
        15'h41FE: data = 12'h508;
        15'h41FF: data = 12'h517;
        15'h4200: data = 12'h529;
        15'h4201: data = 12'h53A;
        15'h4202: data = 12'h553;
        15'h4203: data = 12'h563;
        15'h4204: data = 12'h573;
        15'h4205: data = 12'h58E;
        15'h4206: data = 12'h5A2;
        15'h4207: data = 12'h5BF;
        15'h4208: data = 12'h5CE;
        15'h4209: data = 12'h5EA;
        15'h420A: data = 12'h602;
        15'h420B: data = 12'h61B;
        15'h420C: data = 12'h637;
        15'h420D: data = 12'h64E;
        15'h420E: data = 12'h663;
        15'h420F: data = 12'h67C;
        15'h4210: data = 12'h692;
        15'h4211: data = 12'h6A4;
        15'h4212: data = 12'h6B9;
        15'h4213: data = 12'h6CD;
        15'h4214: data = 12'h6E0;
        15'h4215: data = 12'h6F5;
        15'h4216: data = 12'h70A;
        15'h4217: data = 12'h71E;
        15'h4218: data = 12'h736;
        15'h4219: data = 12'h748;
        15'h421A: data = 12'h75A;
        15'h421B: data = 12'h775;
        15'h421C: data = 12'h78F;
        15'h421D: data = 12'h7A1;
        15'h421E: data = 12'h7BA;
        15'h421F: data = 12'h7D5;
        15'h4220: data = 12'h7F0;
        15'h4221: data = 12'h80A;
        15'h4222: data = 12'h07A;
        15'h4223: data = 12'h08F;
        15'h4224: data = 12'h0A4;
        15'h4225: data = 12'h0B9;
        15'h4226: data = 12'h0D6;
        15'h4227: data = 12'h0EB;
        15'h4228: data = 12'h102;
        15'h4229: data = 12'h112;
        15'h422A: data = 12'h12C;
        15'h422B: data = 12'h145;
        15'h422C: data = 12'h156;
        15'h422D: data = 12'h167;
        15'h422E: data = 12'h17F;
        15'h422F: data = 12'h198;
        15'h4230: data = 12'h1AE;
        15'h4231: data = 12'h1BD;
        15'h4232: data = 12'h1D6;
        15'h4233: data = 12'h1ED;
        15'h4234: data = 12'h204;
        15'h4235: data = 12'h217;
        15'h4236: data = 12'h231;
        15'h4237: data = 12'h248;
        15'h4238: data = 12'h260;
        15'h4239: data = 12'h27B;
        15'h423A: data = 12'h28E;
        15'h423B: data = 12'h2AB;
        15'h423C: data = 12'h2C7;
        15'h423D: data = 12'h2DF;
        15'h423E: data = 12'h2F5;
        15'h423F: data = 12'h30C;
        15'h4240: data = 12'h32A;
        15'h4241: data = 12'h33C;
        15'h4242: data = 12'h352;
        15'h4243: data = 12'h36B;
        15'h4244: data = 12'h37F;
        15'h4245: data = 12'h39F;
        15'h4246: data = 12'h3AE;
        15'h4247: data = 12'h3C2;
        15'h4248: data = 12'h3DA;
        15'h4249: data = 12'h3EF;
        15'h424A: data = 12'h404;
        15'h424B: data = 12'h416;
        15'h424C: data = 12'h428;
        15'h424D: data = 12'h441;
        15'h424E: data = 12'h451;
        15'h424F: data = 12'h465;
        15'h4250: data = 12'h479;
        15'h4251: data = 12'h48F;
        15'h4252: data = 12'h4A4;
        15'h4253: data = 12'h4B4;
        15'h4254: data = 12'h4C3;
        15'h4255: data = 12'h4D9;
        15'h4256: data = 12'h4EE;
        15'h4257: data = 12'h501;
        15'h4258: data = 12'h512;
        15'h4259: data = 12'h527;
        15'h425A: data = 12'h53A;
        15'h425B: data = 12'h54B;
        15'h425C: data = 12'h55C;
        15'h425D: data = 12'h569;
        15'h425E: data = 12'h57F;
        15'h425F: data = 12'h591;
        15'h4260: data = 12'h5A7;
        15'h4261: data = 12'h5BA;
        15'h4262: data = 12'h5C5;
        15'h4263: data = 12'h5D8;
        15'h4264: data = 12'h5EF;
        15'h4265: data = 12'h5FF;
        15'h4266: data = 12'h60F;
        15'h4267: data = 12'h620;
        15'h4268: data = 12'h630;
        15'h4269: data = 12'h644;
        15'h426A: data = 12'h655;
        15'h426B: data = 12'h667;
        15'h426C: data = 12'h676;
        15'h426D: data = 12'h686;
        15'h426E: data = 12'h696;
        15'h426F: data = 12'h6A8;
        15'h4270: data = 12'h6BB;
        15'h4271: data = 12'h6C9;
        15'h4272: data = 12'h6D6;
        15'h4273: data = 12'h6E0;
        15'h4274: data = 12'h6EF;
        15'h4275: data = 12'h700;
        15'h4276: data = 12'h70E;
        15'h4277: data = 12'h716;
        15'h4278: data = 12'h723;
        15'h4279: data = 12'h735;
        15'h427A: data = 12'h73E;
        15'h427B: data = 12'h749;
        15'h427C: data = 12'h74F;
        15'h427D: data = 12'h75E;
        15'h427E: data = 12'h767;
        15'h427F: data = 12'h775;
        15'h4280: data = 12'h77B;
        15'h4281: data = 12'h78D;
        15'h4282: data = 12'h795;
        15'h4283: data = 12'h79C;
        15'h4284: data = 12'h7A3;
        15'h4285: data = 12'h7AD;
        15'h4286: data = 12'h7B3;
        15'h4287: data = 12'h7B9;
        15'h4288: data = 12'h7C4;
        15'h4289: data = 12'h7C9;
        15'h428A: data = 12'h7D1;
        15'h428B: data = 12'h7DC;
        15'h428C: data = 12'h7E0;
        15'h428D: data = 12'h7E9;
        15'h428E: data = 12'h7EC;
        15'h428F: data = 12'h7F2;
        15'h4290: data = 12'h7F7;
        15'h4291: data = 12'h7FB;
        15'h4292: data = 12'h7FB;
        15'h4293: data = 12'h809;
        15'h4294: data = 12'h07C;
        15'h4295: data = 12'h089;
        15'h4296: data = 12'h08F;
        15'h4297: data = 12'h095;
        15'h4298: data = 12'h097;
        15'h4299: data = 12'h0A1;
        15'h429A: data = 12'h0A0;
        15'h429B: data = 12'h0AB;
        15'h429C: data = 12'h0AD;
        15'h429D: data = 12'h0AF;
        15'h429E: data = 12'h0B8;
        15'h429F: data = 12'h0BB;
        15'h42A0: data = 12'h0BD;
        15'h42A1: data = 12'h0BF;
        15'h42A2: data = 12'h0CD;
        15'h42A3: data = 12'h0CD;
        15'h42A4: data = 12'h0D1;
        15'h42A5: data = 12'h0D4;
        15'h42A6: data = 12'h0D5;
        15'h42A7: data = 12'h0D6;
        15'h42A8: data = 12'h0D8;
        15'h42A9: data = 12'h0CC;
        15'h42AA: data = 12'h0CA;
        15'h42AB: data = 12'h0CA;
        15'h42AC: data = 12'h0C6;
        15'h42AD: data = 12'h0BF;
        15'h42AE: data = 12'h0B8;
        15'h42AF: data = 12'h0B2;
        15'h42B0: data = 12'h0AD;
        15'h42B1: data = 12'h0AF;
        15'h42B2: data = 12'h0AA;
        15'h42B3: data = 12'h0AC;
        15'h42B4: data = 12'h0B1;
        15'h42B5: data = 12'h0B3;
        15'h42B6: data = 12'h0AF;
        15'h42B7: data = 12'h0A4;
        15'h42B8: data = 12'h0A2;
        15'h42B9: data = 12'h096;
        15'h42BA: data = 12'h08B;
        15'h42BB: data = 12'h07B;
        15'h42BC: data = 12'h074;
        15'h42BD: data = 12'h077;
        15'h42BE: data = 12'h070;
        15'h42BF: data = 12'h06F;
        15'h42C0: data = 12'h06D;
        15'h42C1: data = 12'h067;
        15'h42C2: data = 12'h060;
        15'h42C3: data = 12'h055;
        15'h42C4: data = 12'h041;
        15'h42C5: data = 12'h034;
        15'h42C6: data = 12'h7B4;
        15'h42C7: data = 12'h7A8;
        15'h42C8: data = 12'h7A6;
        15'h42C9: data = 12'h79D;
        15'h42CA: data = 12'h794;
        15'h42CB: data = 12'h78B;
        15'h42CC: data = 12'h779;
        15'h42CD: data = 12'h768;
        15'h42CE: data = 12'h757;
        15'h42CF: data = 12'h745;
        15'h42D0: data = 12'h736;
        15'h42D1: data = 12'h72F;
        15'h42D2: data = 12'h729;
        15'h42D3: data = 12'h720;
        15'h42D4: data = 12'h714;
        15'h42D5: data = 12'h70B;
        15'h42D6: data = 12'h6FB;
        15'h42D7: data = 12'h6E7;
        15'h42D8: data = 12'h6D6;
        15'h42D9: data = 12'h6C2;
        15'h42DA: data = 12'h6B3;
        15'h42DB: data = 12'h6AA;
        15'h42DC: data = 12'h697;
        15'h42DD: data = 12'h68E;
        15'h42DE: data = 12'h684;
        15'h42DF: data = 12'h677;
        15'h42E0: data = 12'h669;
        15'h42E1: data = 12'h654;
        15'h42E2: data = 12'h645;
        15'h42E3: data = 12'h62F;
        15'h42E4: data = 12'h624;
        15'h42E5: data = 12'h608;
        15'h42E6: data = 12'h5F3;
        15'h42E7: data = 12'h5E1;
        15'h42E8: data = 12'h5CF;
        15'h42E9: data = 12'h5BF;
        15'h42EA: data = 12'h5B6;
        15'h42EB: data = 12'h5A6;
        15'h42EC: data = 12'h596;
        15'h42ED: data = 12'h585;
        15'h42EE: data = 12'h578;
        15'h42EF: data = 12'h569;
        15'h42F0: data = 12'h554;
        15'h42F1: data = 12'h541;
        15'h42F2: data = 12'h529;
        15'h42F3: data = 12'h512;
        15'h42F4: data = 12'h4FF;
        15'h42F5: data = 12'h4EE;
        15'h42F6: data = 12'h4D2;
        15'h42F7: data = 12'h4BA;
        15'h42F8: data = 12'h4A9;
        15'h42F9: data = 12'h491;
        15'h42FA: data = 12'h479;
        15'h42FB: data = 12'h464;
        15'h42FC: data = 12'h451;
        15'h42FD: data = 12'h43E;
        15'h42FE: data = 12'h42A;
        15'h42FF: data = 12'h417;
        15'h4300: data = 12'h404;
        15'h4301: data = 12'h3EE;
        15'h4302: data = 12'h3DD;
        15'h4303: data = 12'h3C7;
        15'h4304: data = 12'h3B4;
        15'h4305: data = 12'h398;
        15'h4306: data = 12'h389;
        15'h4307: data = 12'h373;
        15'h4308: data = 12'h35D;
        15'h4309: data = 12'h348;
        15'h430A: data = 12'h331;
        15'h430B: data = 12'h31C;
        15'h430C: data = 12'h303;
        15'h430D: data = 12'h2F0;
        15'h430E: data = 12'h2DC;
        15'h430F: data = 12'h2C4;
        15'h4310: data = 12'h2A8;
        15'h4311: data = 12'h290;
        15'h4312: data = 12'h280;
        15'h4313: data = 12'h264;
        15'h4314: data = 12'h24C;
        15'h4315: data = 12'h238;
        15'h4316: data = 12'h21B;
        15'h4317: data = 12'h205;
        15'h4318: data = 12'h1EF;
        15'h4319: data = 12'h1D7;
        15'h431A: data = 12'h1BF;
        15'h431B: data = 12'h1AB;
        15'h431C: data = 12'h190;
        15'h431D: data = 12'h17B;
        15'h431E: data = 12'h164;
        15'h431F: data = 12'h14B;
        15'h4320: data = 12'h135;
        15'h4321: data = 12'h118;
        15'h4322: data = 12'h106;
        15'h4323: data = 12'h0EF;
        15'h4324: data = 12'h0D5;
        15'h4325: data = 12'h0B9;
        15'h4326: data = 12'h0A3;
        15'h4327: data = 12'h08C;
        15'h4328: data = 12'h078;
        15'h4329: data = 12'h05E;
        15'h432A: data = 12'h047;
        15'h432B: data = 12'h72A;
        15'h432C: data = 12'h7C8;
        15'h432D: data = 12'h7B3;
        15'h432E: data = 12'h79D;
        15'h432F: data = 12'h789;
        15'h4330: data = 12'h76E;
        15'h4331: data = 12'h756;
        15'h4332: data = 12'h742;
        15'h4333: data = 12'h72F;
        15'h4334: data = 12'h717;
        15'h4335: data = 12'h700;
        15'h4336: data = 12'h6E5;
        15'h4337: data = 12'h6D4;
        15'h4338: data = 12'h6BD;
        15'h4339: data = 12'h6A5;
        15'h433A: data = 12'h68C;
        15'h433B: data = 12'h676;
        15'h433C: data = 12'h65F;
        15'h433D: data = 12'h649;
        15'h433E: data = 12'h630;
        15'h433F: data = 12'h61D;
        15'h4340: data = 12'h605;
        15'h4341: data = 12'h5EC;
        15'h4342: data = 12'h5D6;
        15'h4343: data = 12'h5C0;
        15'h4344: data = 12'h5AC;
        15'h4345: data = 12'h592;
        15'h4346: data = 12'h57B;
        15'h4347: data = 12'h563;
        15'h4348: data = 12'h557;
        15'h4349: data = 12'h543;
        15'h434A: data = 12'h52D;
        15'h434B: data = 12'h51B;
        15'h434C: data = 12'h506;
        15'h434D: data = 12'h4F5;
        15'h434E: data = 12'h4E0;
        15'h434F: data = 12'h4CC;
        15'h4350: data = 12'h4BB;
        15'h4351: data = 12'h4A6;
        15'h4352: data = 12'h497;
        15'h4353: data = 12'h482;
        15'h4354: data = 12'h470;
        15'h4355: data = 12'h462;
        15'h4356: data = 12'h455;
        15'h4357: data = 12'h442;
        15'h4358: data = 12'h42D;
        15'h4359: data = 12'h419;
        15'h435A: data = 12'h40A;
        15'h435B: data = 12'h3F6;
        15'h435C: data = 12'h3E9;
        15'h435D: data = 12'h3CB;
        15'h435E: data = 12'h3BF;
        15'h435F: data = 12'h3A7;
        15'h4360: data = 12'h392;
        15'h4361: data = 12'h387;
        15'h4362: data = 12'h36E;
        15'h4363: data = 12'h35E;
        15'h4364: data = 12'h34D;
        15'h4365: data = 12'h338;
        15'h4366: data = 12'h328;
        15'h4367: data = 12'h31C;
        15'h4368: data = 12'h30D;
        15'h4369: data = 12'h303;
        15'h436A: data = 12'h2F7;
        15'h436B: data = 12'h2EB;
        15'h436C: data = 12'h2DF;
        15'h436D: data = 12'h2DA;
        15'h436E: data = 12'h2CA;
        15'h436F: data = 12'h2BB;
        15'h4370: data = 12'h2AA;
        15'h4371: data = 12'h298;
        15'h4372: data = 12'h292;
        15'h4373: data = 12'h280;
        15'h4374: data = 12'h274;
        15'h4375: data = 12'h261;
        15'h4376: data = 12'h251;
        15'h4377: data = 12'h245;
        15'h4378: data = 12'h239;
        15'h4379: data = 12'h22E;
        15'h437A: data = 12'h223;
        15'h437B: data = 12'h218;
        15'h437C: data = 12'h218;
        15'h437D: data = 12'h213;
        15'h437E: data = 12'h211;
        15'h437F: data = 12'h205;
        15'h4380: data = 12'h1FA;
        15'h4381: data = 12'h1F3;
        15'h4382: data = 12'h1E6;
        15'h4383: data = 12'h1DA;
        15'h4384: data = 12'h1CE;
        15'h4385: data = 12'h1C1;
        15'h4386: data = 12'h1B7;
        15'h4387: data = 12'h1B0;
        15'h4388: data = 12'h1AB;
        15'h4389: data = 12'h1A2;
        15'h438A: data = 12'h19C;
        15'h438B: data = 12'h197;
        15'h438C: data = 12'h19A;
        15'h438D: data = 12'h19A;
        15'h438E: data = 12'h194;
        15'h438F: data = 12'h18D;
        15'h4390: data = 12'h190;
        15'h4391: data = 12'h189;
        15'h4392: data = 12'h185;
        15'h4393: data = 12'h179;
        15'h4394: data = 12'h177;
        15'h4395: data = 12'h16B;
        15'h4396: data = 12'h165;
        15'h4397: data = 12'h163;
        15'h4398: data = 12'h15C;
        15'h4399: data = 12'h15D;
        15'h439A: data = 12'h15E;
        15'h439B: data = 12'h163;
        15'h439C: data = 12'h15E;
        15'h439D: data = 12'h163;
        15'h439E: data = 12'h163;
        15'h439F: data = 12'h168;
        15'h43A0: data = 12'h166;
        15'h43A1: data = 12'h168;
        15'h43A2: data = 12'h167;
        15'h43A3: data = 12'h169;
        15'h43A4: data = 12'h167;
        15'h43A5: data = 12'h166;
        15'h43A6: data = 12'h161;
        15'h43A7: data = 12'h15D;
        15'h43A8: data = 12'h163;
        15'h43A9: data = 12'h161;
        15'h43AA: data = 12'h16E;
        15'h43AB: data = 12'h16E;
        15'h43AC: data = 12'h176;
        15'h43AD: data = 12'h17D;
        15'h43AE: data = 12'h18C;
        15'h43AF: data = 12'h18D;
        15'h43B0: data = 12'h194;
        15'h43B1: data = 12'h198;
        15'h43B2: data = 12'h19C;
        15'h43B3: data = 12'h1A4;
        15'h43B4: data = 12'h1A8;
        15'h43B5: data = 12'h1AD;
        15'h43B6: data = 12'h1A9;
        15'h43B7: data = 12'h1AC;
        15'h43B8: data = 12'h1B1;
        15'h43B9: data = 12'h1B9;
        15'h43BA: data = 12'h1C1;
        15'h43BB: data = 12'h1C8;
        15'h43BC: data = 12'h1D4;
        15'h43BD: data = 12'h1E0;
        15'h43BE: data = 12'h1F1;
        15'h43BF: data = 12'h1FD;
        15'h43C0: data = 12'h207;
        15'h43C1: data = 12'h210;
        15'h43C2: data = 12'h21F;
        15'h43C3: data = 12'h21F;
        15'h43C4: data = 12'h22F;
        15'h43C5: data = 12'h234;
        15'h43C6: data = 12'h23F;
        15'h43C7: data = 12'h243;
        15'h43C8: data = 12'h253;
        15'h43C9: data = 12'h25A;
        15'h43CA: data = 12'h264;
        15'h43CB: data = 12'h26B;
        15'h43CC: data = 12'h27B;
        15'h43CD: data = 12'h28A;
        15'h43CE: data = 12'h293;
        15'h43CF: data = 12'h2A6;
        15'h43D0: data = 12'h2BB;
        15'h43D1: data = 12'h2D1;
        15'h43D2: data = 12'h2DD;
        15'h43D3: data = 12'h2E9;
        15'h43D4: data = 12'h2F9;
        15'h43D5: data = 12'h309;
        15'h43D6: data = 12'h316;
        15'h43D7: data = 12'h326;
        15'h43D8: data = 12'h330;
        15'h43D9: data = 12'h33F;
        15'h43DA: data = 12'h34E;
        15'h43DB: data = 12'h35A;
        15'h43DC: data = 12'h365;
        15'h43DD: data = 12'h373;
        15'h43DE: data = 12'h388;
        15'h43DF: data = 12'h392;
        15'h43E0: data = 12'h3A8;
        15'h43E1: data = 12'h3BA;
        15'h43E2: data = 12'h3CD;
        15'h43E3: data = 12'h3E3;
        15'h43E4: data = 12'h3F5;
        15'h43E5: data = 12'h40C;
        15'h43E6: data = 12'h425;
        15'h43E7: data = 12'h438;
        15'h43E8: data = 12'h44E;
        15'h43E9: data = 12'h45A;
        15'h43EA: data = 12'h46E;
        15'h43EB: data = 12'h481;
        15'h43EC: data = 12'h496;
        15'h43ED: data = 12'h4A8;
        15'h43EE: data = 12'h4B5;
        15'h43EF: data = 12'h4CA;
        15'h43F0: data = 12'h4DD;
        15'h43F1: data = 12'h4F1;
        15'h43F2: data = 12'h500;
        15'h43F3: data = 12'h510;
        15'h43F4: data = 12'h520;
        15'h43F5: data = 12'h539;
        15'h43F6: data = 12'h552;
        15'h43F7: data = 12'h568;
        15'h43F8: data = 12'h577;
        15'h43F9: data = 12'h591;
        15'h43FA: data = 12'h5AB;
        15'h43FB: data = 12'h5C7;
        15'h43FC: data = 12'h5D9;
        15'h43FD: data = 12'h5F1;
        15'h43FE: data = 12'h60B;
        15'h43FF: data = 12'h627;
        15'h4400: data = 12'h63B;
        15'h4401: data = 12'h64F;
        15'h4402: data = 12'h664;
        15'h4403: data = 12'h679;
        15'h4404: data = 12'h690;
        15'h4405: data = 12'h6A1;
        15'h4406: data = 12'h6B1;
        15'h4407: data = 12'h6C7;
        15'h4408: data = 12'h6DB;
        15'h4409: data = 12'h6EC;
        15'h440A: data = 12'h6FF;
        15'h440B: data = 12'h717;
        15'h440C: data = 12'h735;
        15'h440D: data = 12'h743;
        15'h440E: data = 12'h75B;
        15'h440F: data = 12'h777;
        15'h4410: data = 12'h796;
        15'h4411: data = 12'h7A8;
        15'h4412: data = 12'h7C5;
        15'h4413: data = 12'h7E2;
        15'h4414: data = 12'h7FB;
        15'h4415: data = 12'h810;
        15'h4416: data = 12'h07B;
        15'h4417: data = 12'h090;
        15'h4418: data = 12'h0A4;
        15'h4419: data = 12'h0B9;
        15'h441A: data = 12'h0D2;
        15'h441B: data = 12'h0E7;
        15'h441C: data = 12'h0FF;
        15'h441D: data = 12'h10F;
        15'h441E: data = 12'h127;
        15'h441F: data = 12'h13C;
        15'h4420: data = 12'h14F;
        15'h4421: data = 12'h162;
        15'h4422: data = 12'h179;
        15'h4423: data = 12'h192;
        15'h4424: data = 12'h1AB;
        15'h4425: data = 12'h1BC;
        15'h4426: data = 12'h1D8;
        15'h4427: data = 12'h1ED;
        15'h4428: data = 12'h204;
        15'h4429: data = 12'h21A;
        15'h442A: data = 12'h235;
        15'h442B: data = 12'h24E;
        15'h442C: data = 12'h267;
        15'h442D: data = 12'h283;
        15'h442E: data = 12'h297;
        15'h442F: data = 12'h2B3;
        15'h4430: data = 12'h2CA;
        15'h4431: data = 12'h2E5;
        15'h4432: data = 12'h2FD;
        15'h4433: data = 12'h311;
        15'h4434: data = 12'h32B;
        15'h4435: data = 12'h33F;
        15'h4436: data = 12'h352;
        15'h4437: data = 12'h36B;
        15'h4438: data = 12'h380;
        15'h4439: data = 12'h39D;
        15'h443A: data = 12'h3AA;
        15'h443B: data = 12'h3C2;
        15'h443C: data = 12'h3D6;
        15'h443D: data = 12'h3EE;
        15'h443E: data = 12'h3FF;
        15'h443F: data = 12'h411;
        15'h4440: data = 12'h427;
        15'h4441: data = 12'h43D;
        15'h4442: data = 12'h44C;
        15'h4443: data = 12'h45F;
        15'h4444: data = 12'h474;
        15'h4445: data = 12'h48E;
        15'h4446: data = 12'h49E;
        15'h4447: data = 12'h4B1;
        15'h4448: data = 12'h4C3;
        15'h4449: data = 12'h4D6;
        15'h444A: data = 12'h4EA;
        15'h444B: data = 12'h500;
        15'h444C: data = 12'h511;
        15'h444D: data = 12'h52B;
        15'h444E: data = 12'h539;
        15'h444F: data = 12'h54E;
        15'h4450: data = 12'h55B;
        15'h4451: data = 12'h570;
        15'h4452: data = 12'h585;
        15'h4453: data = 12'h595;
        15'h4454: data = 12'h5AE;
        15'h4455: data = 12'h5BF;
        15'h4456: data = 12'h5CE;
        15'h4457: data = 12'h5E0;
        15'h4458: data = 12'h5F6;
        15'h4459: data = 12'h606;
        15'h445A: data = 12'h61A;
        15'h445B: data = 12'h629;
        15'h445C: data = 12'h63C;
        15'h445D: data = 12'h64C;
        15'h445E: data = 12'h65D;
        15'h445F: data = 12'h66B;
        15'h4460: data = 12'h67C;
        15'h4461: data = 12'h689;
        15'h4462: data = 12'h69D;
        15'h4463: data = 12'h6AF;
        15'h4464: data = 12'h6BD;
        15'h4465: data = 12'h6CB;
        15'h4466: data = 12'h6D9;
        15'h4467: data = 12'h6E1;
        15'h4468: data = 12'h6ED;
        15'h4469: data = 12'h700;
        15'h446A: data = 12'h70E;
        15'h446B: data = 12'h714;
        15'h446C: data = 12'h723;
        15'h446D: data = 12'h734;
        15'h446E: data = 12'h73E;
        15'h446F: data = 12'h746;
        15'h4470: data = 12'h753;
        15'h4471: data = 12'h75C;
        15'h4472: data = 12'h765;
        15'h4473: data = 12'h774;
        15'h4474: data = 12'h77B;
        15'h4475: data = 12'h78C;
        15'h4476: data = 12'h790;
        15'h4477: data = 12'h798;
        15'h4478: data = 12'h79D;
        15'h4479: data = 12'h7AA;
        15'h447A: data = 12'h7B1;
        15'h447B: data = 12'h7B3;
        15'h447C: data = 12'h7BC;
        15'h447D: data = 12'h7C6;
        15'h447E: data = 12'h7CD;
        15'h447F: data = 12'h7D4;
        15'h4480: data = 12'h7E2;
        15'h4481: data = 12'h7E4;
        15'h4482: data = 12'h7E7;
        15'h4483: data = 12'h7EE;
        15'h4484: data = 12'h7F5;
        15'h4485: data = 12'h7FC;
        15'h4486: data = 12'h7FE;
        15'h4487: data = 12'h805;
        15'h4488: data = 12'h4CD;
        15'h4489: data = 12'h084;
        15'h448A: data = 12'h08E;
        15'h448B: data = 12'h093;
        15'h448C: data = 12'h098;
        15'h448D: data = 12'h09F;
        15'h448E: data = 12'h0A1;
        15'h448F: data = 12'h0AC;
        15'h4490: data = 12'h0AC;
        15'h4491: data = 12'h0AF;
        15'h4492: data = 12'h0BB;
        15'h4493: data = 12'h0BD;
        15'h4494: data = 12'h0C2;
        15'h4495: data = 12'h0C6;
        15'h4496: data = 12'h0D1;
        15'h4497: data = 12'h0D7;
        15'h4498: data = 12'h0D4;
        15'h4499: data = 12'h0D8;
        15'h449A: data = 12'h0D7;
        15'h449B: data = 12'h0D5;
        15'h449C: data = 12'h0D3;
        15'h449D: data = 12'h0CA;
        15'h449E: data = 12'h0C9;
        15'h449F: data = 12'h0C7;
        15'h44A0: data = 12'h0C5;
        15'h44A1: data = 12'h0BC;
        15'h44A2: data = 12'h0B4;
        15'h44A3: data = 12'h0B4;
        15'h44A4: data = 12'h0AF;
        15'h44A5: data = 12'h0B3;
        15'h44A6: data = 12'h0B1;
        15'h44A7: data = 12'h0B6;
        15'h44A8: data = 12'h0B8;
        15'h44A9: data = 12'h0B8;
        15'h44AA: data = 12'h0AF;
        15'h44AB: data = 12'h0A5;
        15'h44AC: data = 12'h0A1;
        15'h44AD: data = 12'h096;
        15'h44AE: data = 12'h08A;
        15'h44AF: data = 12'h07E;
        15'h44B0: data = 12'h078;
        15'h44B1: data = 12'h077;
        15'h44B2: data = 12'h078;
        15'h44B3: data = 12'h075;
        15'h44B4: data = 12'h06D;
        15'h44B5: data = 12'h068;
        15'h44B6: data = 12'h061;
        15'h44B7: data = 12'h050;
        15'h44B8: data = 12'h03C;
        15'h44B9: data = 12'h030;
        15'h44BA: data = 12'h7B6;
        15'h44BB: data = 12'h7AA;
        15'h44BC: data = 12'h7AC;
        15'h44BD: data = 12'h7A1;
        15'h44BE: data = 12'h798;
        15'h44BF: data = 12'h789;
        15'h44C0: data = 12'h77B;
        15'h44C1: data = 12'h768;
        15'h44C2: data = 12'h753;
        15'h44C3: data = 12'h741;
        15'h44C4: data = 12'h734;
        15'h44C5: data = 12'h730;
        15'h44C6: data = 12'h72D;
        15'h44C7: data = 12'h723;
        15'h44C8: data = 12'h717;
        15'h44C9: data = 12'h70B;
        15'h44CA: data = 12'h6FA;
        15'h44CB: data = 12'h6E5;
        15'h44CC: data = 12'h6D1;
        15'h44CD: data = 12'h6C2;
        15'h44CE: data = 12'h6B1;
        15'h44CF: data = 12'h6A4;
        15'h44D0: data = 12'h696;
        15'h44D1: data = 12'h68E;
        15'h44D2: data = 12'h685;
        15'h44D3: data = 12'h675;
        15'h44D4: data = 12'h669;
        15'h44D5: data = 12'h658;
        15'h44D6: data = 12'h642;
        15'h44D7: data = 12'h62D;
        15'h44D8: data = 12'h622;
        15'h44D9: data = 12'h607;
        15'h44DA: data = 12'h5F6;
        15'h44DB: data = 12'h5E5;
        15'h44DC: data = 12'h5D2;
        15'h44DD: data = 12'h5C5;
        15'h44DE: data = 12'h5BB;
        15'h44DF: data = 12'h5A9;
        15'h44E0: data = 12'h599;
        15'h44E1: data = 12'h586;
        15'h44E2: data = 12'h576;
        15'h44E3: data = 12'h567;
        15'h44E4: data = 12'h556;
        15'h44E5: data = 12'h53F;
        15'h44E6: data = 12'h52A;
        15'h44E7: data = 12'h513;
        15'h44E8: data = 12'h4FC;
        15'h44E9: data = 12'h4E8;
        15'h44EA: data = 12'h4CE;
        15'h44EB: data = 12'h4B5;
        15'h44EC: data = 12'h4A4;
        15'h44ED: data = 12'h490;
        15'h44EE: data = 12'h47B;
        15'h44EF: data = 12'h465;
        15'h44F0: data = 12'h451;
        15'h44F1: data = 12'h442;
        15'h44F2: data = 12'h42D;
        15'h44F3: data = 12'h41B;
        15'h44F4: data = 12'h408;
        15'h44F5: data = 12'h3F3;
        15'h44F6: data = 12'h3DB;
        15'h44F7: data = 12'h3CA;
        15'h44F8: data = 12'h3B3;
        15'h44F9: data = 12'h39D;
        15'h44FA: data = 12'h38F;
        15'h44FB: data = 12'h375;
        15'h44FC: data = 12'h35E;
        15'h44FD: data = 12'h348;
        15'h44FE: data = 12'h332;
        15'h44FF: data = 12'h31D;
        15'h4500: data = 12'h307;
        15'h4501: data = 12'h2F0;
        15'h4502: data = 12'h2DB;
        15'h4503: data = 12'h2C5;
        15'h4504: data = 12'h2A7;
        15'h4505: data = 12'h295;
        15'h4506: data = 12'h280;
        15'h4507: data = 12'h264;
        15'h4508: data = 12'h24A;
        15'h4509: data = 12'h234;
        15'h450A: data = 12'h21E;
        15'h450B: data = 12'h203;
        15'h450C: data = 12'h1EE;
        15'h450D: data = 12'h1D5;
        15'h450E: data = 12'h1C0;
        15'h450F: data = 12'h1A5;
        15'h4510: data = 12'h18F;
        15'h4511: data = 12'h179;
        15'h4512: data = 12'h162;
        15'h4513: data = 12'h14A;
        15'h4514: data = 12'h131;
        15'h4515: data = 12'h117;
        15'h4516: data = 12'h103;
        15'h4517: data = 12'h0F0;
        15'h4518: data = 12'h0D4;
        15'h4519: data = 12'h0BC;
        15'h451A: data = 12'h0A4;
        15'h451B: data = 12'h08C;
        15'h451C: data = 12'h077;
        15'h451D: data = 12'h05D;
        15'h451E: data = 12'h046;
        15'h451F: data = 12'h75E;
        15'h4520: data = 12'h7C7;
        15'h4521: data = 12'h7B2;
        15'h4522: data = 12'h79D;
        15'h4523: data = 12'h786;
        15'h4524: data = 12'h76F;
        15'h4525: data = 12'h754;
        15'h4526: data = 12'h741;
        15'h4527: data = 12'h72E;
        15'h4528: data = 12'h718;
        15'h4529: data = 12'h6FD;
        15'h452A: data = 12'h6E0;
        15'h452B: data = 12'h6CD;
        15'h452C: data = 12'h6BB;
        15'h452D: data = 12'h6A3;
        15'h452E: data = 12'h686;
        15'h452F: data = 12'h675;
        15'h4530: data = 12'h65B;
        15'h4531: data = 12'h64A;
        15'h4532: data = 12'h633;
        15'h4533: data = 12'h61B;
        15'h4534: data = 12'h604;
        15'h4535: data = 12'h5E9;
        15'h4536: data = 12'h5D5;
        15'h4537: data = 12'h5C2;
        15'h4538: data = 12'h5AB;
        15'h4539: data = 12'h593;
        15'h453A: data = 12'h57E;
        15'h453B: data = 12'h56A;
        15'h453C: data = 12'h559;
        15'h453D: data = 12'h540;
        15'h453E: data = 12'h52D;
        15'h453F: data = 12'h51C;
        15'h4540: data = 12'h50C;
        15'h4541: data = 12'h4F7;
        15'h4542: data = 12'h4E2;
        15'h4543: data = 12'h4CF;
        15'h4544: data = 12'h4BC;
        15'h4545: data = 12'h4AC;
        15'h4546: data = 12'h49F;
        15'h4547: data = 12'h48B;
        15'h4548: data = 12'h477;
        15'h4549: data = 12'h465;
        15'h454A: data = 12'h458;
        15'h454B: data = 12'h441;
        15'h454C: data = 12'h432;
        15'h454D: data = 12'h419;
        15'h454E: data = 12'h406;
        15'h454F: data = 12'h3F8;
        15'h4550: data = 12'h3E3;
        15'h4551: data = 12'h3CE;
        15'h4552: data = 12'h3BD;
        15'h4553: data = 12'h3A5;
        15'h4554: data = 12'h391;
        15'h4555: data = 12'h385;
        15'h4556: data = 12'h36F;
        15'h4557: data = 12'h35C;
        15'h4558: data = 12'h34C;
        15'h4559: data = 12'h33F;
        15'h455A: data = 12'h32D;
        15'h455B: data = 12'h320;
        15'h455C: data = 12'h314;
        15'h455D: data = 12'h307;
        15'h455E: data = 12'h2FA;
        15'h455F: data = 12'h2F0;
        15'h4560: data = 12'h2E6;
        15'h4561: data = 12'h2DA;
        15'h4562: data = 12'h2CC;
        15'h4563: data = 12'h2BF;
        15'h4564: data = 12'h2AC;
        15'h4565: data = 12'h29C;
        15'h4566: data = 12'h28F;
        15'h4567: data = 12'h27C;
        15'h4568: data = 12'h26F;
        15'h4569: data = 12'h25E;
        15'h456A: data = 12'h255;
        15'h456B: data = 12'h244;
        15'h456C: data = 12'h23B;
        15'h456D: data = 12'h231;
        15'h456E: data = 12'h224;
        15'h456F: data = 12'h21F;
        15'h4570: data = 12'h21B;
        15'h4571: data = 12'h216;
        15'h4572: data = 12'h20C;
        15'h4573: data = 12'h200;
        15'h4574: data = 12'h1FA;
        15'h4575: data = 12'h1EF;
        15'h4576: data = 12'h1E6;
        15'h4577: data = 12'h1DA;
        15'h4578: data = 12'h1CA;
        15'h4579: data = 12'h1C0;
        15'h457A: data = 12'h1B1;
        15'h457B: data = 12'h1B2;
        15'h457C: data = 12'h1AB;
        15'h457D: data = 12'h1A5;
        15'h457E: data = 12'h19D;
        15'h457F: data = 12'h19B;
        15'h4580: data = 12'h19C;
        15'h4581: data = 12'h19D;
        15'h4582: data = 12'h195;
        15'h4583: data = 12'h18F;
        15'h4584: data = 12'h18F;
        15'h4585: data = 12'h186;
        15'h4586: data = 12'h184;
        15'h4587: data = 12'h177;
        15'h4588: data = 12'h175;
        15'h4589: data = 12'h169;
        15'h458A: data = 12'h168;
        15'h458B: data = 12'h167;
        15'h458C: data = 12'h15C;
        15'h458D: data = 12'h160;
        15'h458E: data = 12'h163;
        15'h458F: data = 12'h167;
        15'h4590: data = 12'h163;
        15'h4591: data = 12'h165;
        15'h4592: data = 12'h169;
        15'h4593: data = 12'h167;
        15'h4594: data = 12'h166;
        15'h4595: data = 12'h165;
        15'h4596: data = 12'h167;
        15'h4597: data = 12'h16A;
        15'h4598: data = 12'h164;
        15'h4599: data = 12'h161;
        15'h459A: data = 12'h161;
        15'h459B: data = 12'h15F;
        15'h459C: data = 12'h163;
        15'h459D: data = 12'h167;
        15'h459E: data = 12'h171;
        15'h459F: data = 12'h175;
        15'h45A0: data = 12'h17F;
        15'h45A1: data = 12'h186;
        15'h45A2: data = 12'h18F;
        15'h45A3: data = 12'h18D;
        15'h45A4: data = 12'h196;
        15'h45A5: data = 12'h198;
        15'h45A6: data = 12'h199;
        15'h45A7: data = 12'h1A0;
        15'h45A8: data = 12'h1A7;
        15'h45A9: data = 12'h1A9;
        15'h45AA: data = 12'h1A9;
        15'h45AB: data = 12'h1AB;
        15'h45AC: data = 12'h1AF;
        15'h45AD: data = 12'h1BA;
        15'h45AE: data = 12'h1C4;
        15'h45AF: data = 12'h1CA;
        15'h45B0: data = 12'h1D8;
        15'h45B1: data = 12'h1E5;
        15'h45B2: data = 12'h1F4;
        15'h45B3: data = 12'h202;
        15'h45B4: data = 12'h209;
        15'h45B5: data = 12'h212;
        15'h45B6: data = 12'h222;
        15'h45B7: data = 12'h21F;
        15'h45B8: data = 12'h231;
        15'h45B9: data = 12'h233;
        15'h45BA: data = 12'h241;
        15'h45BB: data = 12'h241;
        15'h45BC: data = 12'h24F;
        15'h45BD: data = 12'h25A;
        15'h45BE: data = 12'h262;
        15'h45BF: data = 12'h26D;
        15'h45C0: data = 12'h279;
        15'h45C1: data = 12'h28C;
        15'h45C2: data = 12'h298;
        15'h45C3: data = 12'h2AC;
        15'h45C4: data = 12'h2BE;
        15'h45C5: data = 12'h2CF;
        15'h45C6: data = 12'h2E1;
        15'h45C7: data = 12'h2EB;
        15'h45C8: data = 12'h2FA;
        15'h45C9: data = 12'h309;
        15'h45CA: data = 12'h318;
        15'h45CB: data = 12'h325;
        15'h45CC: data = 12'h333;
        15'h45CD: data = 12'h33E;
        15'h45CE: data = 12'h349;
        15'h45CF: data = 12'h357;
        15'h45D0: data = 12'h368;
        15'h45D1: data = 12'h373;
        15'h45D2: data = 12'h389;
        15'h45D3: data = 12'h395;
        15'h45D4: data = 12'h3AA;
        15'h45D5: data = 12'h3B8;
        15'h45D6: data = 12'h3CF;
        15'h45D7: data = 12'h3E5;
        15'h45D8: data = 12'h3FA;
        15'h45D9: data = 12'h40D;
        15'h45DA: data = 12'h425;
        15'h45DB: data = 12'h436;
        15'h45DC: data = 12'h44B;
        15'h45DD: data = 12'h45C;
        15'h45DE: data = 12'h46E;
        15'h45DF: data = 12'h482;
        15'h45E0: data = 12'h493;
        15'h45E1: data = 12'h4A5;
        15'h45E2: data = 12'h4B2;
        15'h45E3: data = 12'h4C4;
        15'h45E4: data = 12'h4D6;
        15'h45E5: data = 12'h4E8;
        15'h45E6: data = 12'h4FC;
        15'h45E7: data = 12'h512;
        15'h45E8: data = 12'h524;
        15'h45E9: data = 12'h538;
        15'h45EA: data = 12'h553;
        15'h45EB: data = 12'h568;
        15'h45EC: data = 12'h57E;
        15'h45ED: data = 12'h596;
        15'h45EE: data = 12'h5AF;
        15'h45EF: data = 12'h5C8;
        15'h45F0: data = 12'h5D8;
        15'h45F1: data = 12'h5F5;
        15'h45F2: data = 12'h60C;
        15'h45F3: data = 12'h620;
        15'h45F4: data = 12'h637;
        15'h45F5: data = 12'h64B;
        15'h45F6: data = 12'h661;
        15'h45F7: data = 12'h678;
        15'h45F8: data = 12'h689;
        15'h45F9: data = 12'h69B;
        15'h45FA: data = 12'h6AC;
        15'h45FB: data = 12'h6C6;
        15'h45FC: data = 12'h6D5;
        15'h45FD: data = 12'h6EB;
        15'h45FE: data = 12'h6FD;
        15'h45FF: data = 12'h719;
        15'h4600: data = 12'h736;
        15'h4601: data = 12'h744;
        15'h4602: data = 12'h75F;
        15'h4603: data = 12'h77C;
        15'h4604: data = 12'h79A;
        15'h4605: data = 12'h7AD;
        15'h4606: data = 12'h7C9;
        15'h4607: data = 12'h7E5;
        15'h4608: data = 12'h7FB;
        15'h4609: data = 12'h80F;
        15'h460A: data = 12'h07D;
        15'h460B: data = 12'h092;
        15'h460C: data = 12'h0A5;
        15'h460D: data = 12'h0BA;
        15'h460E: data = 12'h0CE;
        15'h460F: data = 12'h0E6;
        15'h4610: data = 12'h0F8;
        15'h4611: data = 12'h10A;
        15'h4612: data = 12'h122;
        15'h4613: data = 12'h13B;
        15'h4614: data = 12'h14A;
        15'h4615: data = 12'h15F;
        15'h4616: data = 12'h177;
        15'h4617: data = 12'h191;
        15'h4618: data = 12'h1A8;
        15'h4619: data = 12'h1B9;
        15'h461A: data = 12'h1D7;
        15'h461B: data = 12'h1F1;
        15'h461C: data = 12'h208;
        15'h461D: data = 12'h221;
        15'h461E: data = 12'h23B;
        15'h461F: data = 12'h256;
        15'h4620: data = 12'h26E;
        15'h4621: data = 12'h286;
        15'h4622: data = 12'h29C;
        15'h4623: data = 12'h2B6;
        15'h4624: data = 12'h2CF;
        15'h4625: data = 12'h2E8;
        15'h4626: data = 12'h2FF;
        15'h4627: data = 12'h313;
        15'h4628: data = 12'h327;
        15'h4629: data = 12'h340;
        15'h462A: data = 12'h350;
        15'h462B: data = 12'h36D;
        15'h462C: data = 12'h381;
        15'h462D: data = 12'h396;
        15'h462E: data = 12'h3A8;
        15'h462F: data = 12'h3C0;
        15'h4630: data = 12'h3D2;
        15'h4631: data = 12'h3E5;
        15'h4632: data = 12'h3F5;
        15'h4633: data = 12'h40B;
        15'h4634: data = 12'h41F;
        15'h4635: data = 12'h436;
        15'h4636: data = 12'h448;
        15'h4637: data = 12'h459;
        15'h4638: data = 12'h46E;
        15'h4639: data = 12'h48A;
        15'h463A: data = 12'h4A1;
        15'h463B: data = 12'h4AE;
        15'h463C: data = 12'h4C3;
        15'h463D: data = 12'h4D4;
        15'h463E: data = 12'h4EC;
        15'h463F: data = 12'h505;
        15'h4640: data = 12'h513;
        15'h4641: data = 12'h529;
        15'h4642: data = 12'h53C;
        15'h4643: data = 12'h54F;
        15'h4644: data = 12'h560;
        15'h4645: data = 12'h575;
        15'h4646: data = 12'h589;
        15'h4647: data = 12'h59A;
        15'h4648: data = 12'h5B6;
        15'h4649: data = 12'h5C4;
        15'h464A: data = 12'h5D6;
        15'h464B: data = 12'h5E3;
        15'h464C: data = 12'h5FC;
        15'h464D: data = 12'h60B;
        15'h464E: data = 12'h61B;
        15'h464F: data = 12'h62B;
        15'h4650: data = 12'h63C;
        15'h4651: data = 12'h64F;
        15'h4652: data = 12'h65F;
        15'h4653: data = 12'h66E;
        15'h4654: data = 12'h680;
        15'h4655: data = 12'h68E;
        15'h4656: data = 12'h69B;
        15'h4657: data = 12'h6AB;
        15'h4658: data = 12'h6BB;
        15'h4659: data = 12'h6C6;
        15'h465A: data = 12'h6D8;
        15'h465B: data = 12'h6DE;
        15'h465C: data = 12'h6EE;
        15'h465D: data = 12'h6FD;
        15'h465E: data = 12'h709;
        15'h465F: data = 12'h714;
        15'h4660: data = 12'h724;
        15'h4661: data = 12'h733;
        15'h4662: data = 12'h739;
        15'h4663: data = 12'h746;
        15'h4664: data = 12'h74D;
        15'h4665: data = 12'h75A;
        15'h4666: data = 12'h762;
        15'h4667: data = 12'h76C;
        15'h4668: data = 12'h774;
        15'h4669: data = 12'h782;
        15'h466A: data = 12'h788;
        15'h466B: data = 12'h792;
        15'h466C: data = 12'h796;
        15'h466D: data = 12'h7A6;
        15'h466E: data = 12'h7A9;
        15'h466F: data = 12'h7B2;
        15'h4670: data = 12'h7B9;
        15'h4671: data = 12'h7BF;
        15'h4672: data = 12'h7C7;
        15'h4673: data = 12'h7D0;
        15'h4674: data = 12'h7DA;
        15'h4675: data = 12'h7DF;
        15'h4676: data = 12'h7E5;
        15'h4677: data = 12'h7EB;
        15'h4678: data = 12'h7F5;
        15'h4679: data = 12'h7FB;
        15'h467A: data = 12'h7F9;
        15'h467B: data = 12'h500;
        15'h467C: data = 12'h085;
        15'h467D: data = 12'h087;
        15'h467E: data = 12'h093;
        15'h467F: data = 12'h099;
        15'h4680: data = 12'h098;
        15'h4681: data = 12'h0A5;
        15'h4682: data = 12'h0AB;
        15'h4683: data = 12'h0B1;
        15'h4684: data = 12'h0B6;
        15'h4685: data = 12'h0B8;
        15'h4686: data = 12'h0C5;
        15'h4687: data = 12'h0C6;
        15'h4688: data = 12'h0C8;
        15'h4689: data = 12'h0CC;
        15'h468A: data = 12'h0D2;
        15'h468B: data = 12'h0D5;
        15'h468C: data = 12'h0D5;
        15'h468D: data = 12'h0D6;
        15'h468E: data = 12'h0D2;
        15'h468F: data = 12'h0D1;
        15'h4690: data = 12'h0CF;
        15'h4691: data = 12'h0C3;
        15'h4692: data = 12'h0C1;
        15'h4693: data = 12'h0BD;
        15'h4694: data = 12'h0BC;
        15'h4695: data = 12'h0B6;
        15'h4696: data = 12'h0B5;
        15'h4697: data = 12'h0B8;
        15'h4698: data = 12'h0B6;
        15'h4699: data = 12'h0BA;
        15'h469A: data = 12'h0B1;
        15'h469B: data = 12'h0B9;
        15'h469C: data = 12'h0B7;
        15'h469D: data = 12'h0B4;
        15'h469E: data = 12'h0A9;
        15'h469F: data = 12'h09E;
        15'h46A0: data = 12'h097;
        15'h46A1: data = 12'h089;
        15'h46A2: data = 12'h082;
        15'h46A3: data = 12'h07C;
        15'h46A4: data = 12'h078;
        15'h46A5: data = 12'h080;
        15'h46A6: data = 12'h07B;
        15'h46A7: data = 12'h074;
        15'h46A8: data = 12'h06F;
        15'h46A9: data = 12'h063;
        15'h46AA: data = 12'h056;
        15'h46AB: data = 12'h043;
        15'h46AC: data = 12'h036;
        15'h46AD: data = 12'h020;
        15'h46AE: data = 12'h7B5;
        15'h46AF: data = 12'h7B4;
        15'h46B0: data = 12'h7B1;
        15'h46B1: data = 12'h7A2;
        15'h46B2: data = 12'h796;
        15'h46B3: data = 12'h785;
        default: data = 12'h000;
    endcase
end

endmodule

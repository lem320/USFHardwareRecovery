module rom_test2 (
    input [14:0] address,
    output reg [11:0] data
);

always @(*) begin
    case (address)
        15'h0000: data = 12'h3E4;
        15'h0001: data = 12'h32A;
        15'h0002: data = 12'h268;
        15'h0003: data = 12'h196;
        15'h0004: data = 12'h0BC;
        15'h0005: data = 12'h799;
        15'h0006: data = 12'h6A6;
        15'h0007: data = 12'h5A2;
        15'h0008: data = 12'h49C;
        15'h0009: data = 12'h37B;
        15'h000A: data = 12'h265;
        15'h000B: data = 12'h144;
        15'h000C: data = 12'h021;
        15'h000D: data = 12'h6B4;
        15'h000E: data = 12'h586;
        15'h000F: data = 12'h473;
        15'h0010: data = 12'h353;
        15'h0011: data = 12'h241;
        15'h0012: data = 12'h12D;
        15'h0013: data = 12'h031;
        15'h0014: data = 12'h708;
        15'h0015: data = 12'h620;
        15'h0016: data = 12'h53C;
        15'h0017: data = 12'h470;
        15'h0018: data = 12'h39D;
        15'h0019: data = 12'h2E2;
        15'h001A: data = 12'h233;
        15'h001B: data = 12'h1A2;
        15'h001C: data = 12'h10B;
        15'h001D: data = 12'h50D;
        15'h001E: data = 12'h5F7;
        15'h001F: data = 12'h783;
        15'h0020: data = 12'h782;
        15'h0021: data = 12'h764;
        15'h0022: data = 12'h786;
        15'h0023: data = 12'h7A1;
        15'h0024: data = 12'h7E1;
        15'h0025: data = 12'h092;
        15'h0026: data = 12'h0F6;
        15'h0027: data = 12'h16A;
        15'h0028: data = 12'h1FF;
        15'h0029: data = 12'h2A7;
        15'h002A: data = 12'h35D;
        15'h002B: data = 12'h432;
        15'h002C: data = 12'h506;
        15'h002D: data = 12'h5E5;
        15'h002E: data = 12'h6CE;
        15'h002F: data = 12'h7C5;
        15'h0030: data = 12'h0F1;
        15'h0031: data = 12'h1F9;
        15'h0032: data = 12'h2FF;
        15'h0033: data = 12'h422;
        15'h0034: data = 12'h535;
        15'h0035: data = 12'h664;
        15'h0036: data = 12'h78E;
        15'h0037: data = 12'h0EE;
        15'h0038: data = 12'h218;
        15'h0039: data = 12'h331;
        15'h003A: data = 12'h446;
        15'h003B: data = 12'h553;
        15'h003C: data = 12'h50D;
        15'h003D: data = 12'h74D;
        15'h003E: data = 12'h29D;
        15'h003F: data = 12'h160;
        15'h0040: data = 12'h238;
        15'h0041: data = 12'h302;
        15'h0042: data = 12'h3BA;
        15'h0043: data = 12'h45F;
        15'h0044: data = 12'h4EB;
        15'h0045: data = 12'h55D;
        15'h0046: data = 12'h5CA;
        15'h0047: data = 12'h609;
        15'h0048: data = 12'h649;
        15'h0049: data = 12'h671;
        15'h004A: data = 12'h686;
        15'h004B: data = 12'h68A;
        15'h004C: data = 12'h671;
        15'h004D: data = 12'h64A;
        15'h004E: data = 12'h5FA;
        15'h004F: data = 12'h5AA;
        15'h0050: data = 12'h53B;
        15'h0051: data = 12'h4B2;
        15'h0052: data = 12'h410;
        15'h0053: data = 12'h362;
        15'h0054: data = 12'h2A6;
        15'h0055: data = 12'h1DC;
        15'h0056: data = 12'h106;
        15'h0057: data = 12'h05B;
        15'h0058: data = 12'h6F5;
        15'h0059: data = 12'h5FE;
        15'h005A: data = 12'h4F5;
        15'h005B: data = 12'h50D;
        15'h005C: data = 12'h2C2;
        15'h005D: data = 12'h1A9;
        15'h005E: data = 12'h086;
        15'h005F: data = 12'h705;
        15'h0060: data = 12'h5F0;
        15'h0061: data = 12'h4D6;
        15'h0062: data = 12'h3B2;
        15'h0063: data = 12'h2A2;
        15'h0064: data = 12'h18D;
        15'h0065: data = 12'h090;
        15'h0066: data = 12'h75A;
        15'h0067: data = 12'h675;
        15'h0068: data = 12'h583;
        15'h0069: data = 12'h4B2;
        15'h006A: data = 12'h3DF;
        15'h006B: data = 12'h31E;
        15'h006C: data = 12'h274;
        15'h006D: data = 12'h1CD;
        15'h006E: data = 12'h13E;
        15'h006F: data = 12'h0D5;
        15'h0070: data = 12'h076;
        15'h0071: data = 12'h033;
        15'h0072: data = 12'h7A4;
        15'h0073: data = 12'h787;
        15'h0074: data = 12'h764;
        15'h0075: data = 12'h784;
        15'h0076: data = 12'h7A2;
        15'h0077: data = 12'h7D7;
        15'h0078: data = 12'h672;
        15'h0079: data = 12'h0D6;
        15'h007A: data = 12'h50D;
        15'h007B: data = 12'h1CB;
        15'h007C: data = 12'h270;
        15'h007D: data = 12'h328;
        15'h007E: data = 12'h3E5;
        15'h007F: data = 12'h4BC;
        15'h0080: data = 12'h591;
        15'h0081: data = 12'h680;
        15'h0082: data = 12'h76F;
        15'h0083: data = 12'h1C2;
        15'h0084: data = 12'h19B;
        15'h0085: data = 12'h2B5;
        15'h0086: data = 12'h3C5;
        15'h0087: data = 12'h4E9;
        15'h0088: data = 12'h601;
        15'h0089: data = 12'h722;
        15'h008A: data = 12'h7B8;
        15'h008B: data = 12'h1BB;
        15'h008C: data = 12'h2D6;
        15'h008D: data = 12'h3F6;
        15'h008E: data = 12'h503;
        15'h008F: data = 12'h5FC;
        15'h0090: data = 12'h6F8;
        15'h0091: data = 12'h7F0;
        15'h0092: data = 12'h111;
        15'h0093: data = 12'h1EE;
        15'h0094: data = 12'h2BB;
        15'h0095: data = 12'h37A;
        15'h0096: data = 12'h425;
        15'h0097: data = 12'h4BF;
        15'h0098: data = 12'h53E;
        15'h0099: data = 12'h50D;
        15'h009A: data = 12'h5EE;
        15'h009B: data = 12'h63B;
        15'h009C: data = 12'h667;
        15'h009D: data = 12'h688;
        15'h009E: data = 12'h686;
        15'h009F: data = 12'h679;
        15'h00A0: data = 12'h654;
        15'h00A1: data = 12'h616;
        15'h00A2: data = 12'h5CB;
        15'h00A3: data = 12'h558;
        15'h00A4: data = 12'h4DF;
        15'h00A5: data = 12'h453;
        15'h00A6: data = 12'h3A5;
        15'h00A7: data = 12'h2EA;
        15'h00A8: data = 12'h220;
        15'h00A9: data = 12'h150;
        15'h00AA: data = 12'h06B;
        15'h00AB: data = 12'h73C;
        15'h00AC: data = 12'h648;
        15'h00AD: data = 12'h54C;
        15'h00AE: data = 12'h43D;
        15'h00AF: data = 12'h32F;
        15'h00B0: data = 12'h211;
        15'h00B1: data = 12'h0EF;
        15'h00B2: data = 12'h76D;
        15'h00B3: data = 12'h64D;
        15'h00B4: data = 12'h52F;
        15'h00B5: data = 12'h416;
        15'h00B6: data = 12'h2F5;
        15'h00B7: data = 12'h1E2;
        15'h00B8: data = 12'h50D;
        15'h00B9: data = 12'h799;
        15'h00BA: data = 12'h6BF;
        15'h00BB: data = 12'h5D5;
        15'h00BC: data = 12'h4FA;
        15'h00BD: data = 12'h421;
        15'h00BE: data = 12'h35B;
        15'h00BF: data = 12'h2AB;
        15'h00C0: data = 12'h200;
        15'h00C1: data = 12'h170;
        15'h00C2: data = 12'h0F7;
        15'h00C3: data = 12'h098;
        15'h00C4: data = 12'h03D;
        15'h00C5: data = 12'h799;
        15'h00C6: data = 12'h77F;
        15'h00C7: data = 12'h760;
        15'h00C8: data = 12'h782;
        15'h00C9: data = 12'h781;
        15'h00CA: data = 12'h7C2;
        15'h00CB: data = 12'h803;
        15'h00CC: data = 12'h0C0;
        15'h00CD: data = 12'h116;
        15'h00CE: data = 12'h1A3;
        15'h00CF: data = 12'h235;
        15'h00D0: data = 12'h2E0;
        15'h00D1: data = 12'h39D;
        15'h00D2: data = 12'h470;
        15'h00D3: data = 12'h544;
        15'h00D4: data = 12'h632;
        15'h00D5: data = 12'h722;
        15'h00D6: data = 12'h81C;
        15'h00D7: data = 12'h50D;
        15'h00D8: data = 12'h257;
        15'h00D9: data = 12'h36A;
        15'h00DA: data = 12'h480;
        15'h00DB: data = 12'h599;
        15'h00DC: data = 12'h6C2;
        15'h00DD: data = 12'h7E2;
        15'h00DE: data = 12'h154;
        15'h00DF: data = 12'h27B;
        15'h00E0: data = 12'h393;
        15'h00E1: data = 12'h4A8;
        15'h00E2: data = 12'h5AB;
        15'h00E3: data = 12'h6B3;
        15'h00E4: data = 12'h799;
        15'h00E5: data = 12'h0CB;
        15'h00E6: data = 12'h1A3;
        15'h00E7: data = 12'h275;
        15'h00E8: data = 12'h338;
        15'h00E9: data = 12'h3F4;
        15'h00EA: data = 12'h492;
        15'h00EB: data = 12'h51E;
        15'h00EC: data = 12'h589;
        15'h00ED: data = 12'h5EF;
        15'h00EE: data = 12'h632;
        15'h00EF: data = 12'h669;
        15'h00F0: data = 12'h68A;
        15'h00F1: data = 12'h684;
        15'h00F2: data = 12'h685;
        15'h00F3: data = 12'h668;
        15'h00F4: data = 12'h631;
        15'h00F5: data = 12'h5EB;
        15'h00F6: data = 12'h50D;
        15'h00F7: data = 12'h512;
        15'h00F8: data = 12'h484;
        15'h00F9: data = 12'h3E7;
        15'h00FA: data = 12'h334;
        15'h00FB: data = 12'h26F;
        15'h00FC: data = 12'h194;
        15'h00FD: data = 12'h0BB;
        15'h00FE: data = 12'h790;
        15'h00FF: data = 12'h69D;
        15'h0100: data = 12'h598;
        15'h0101: data = 12'h497;
        15'h0102: data = 12'h37A;
        15'h0103: data = 12'h267;
        15'h0104: data = 12'h14C;
        15'h0105: data = 12'h02D;
        15'h0106: data = 12'h6C6;
        15'h0107: data = 12'h594;
        15'h0108: data = 12'h47A;
        15'h0109: data = 12'h359;
        15'h010A: data = 12'h23C;
        15'h010B: data = 12'h12A;
        15'h010C: data = 12'h02B;
        15'h010D: data = 12'h70B;
        15'h010E: data = 12'h615;
        15'h010F: data = 12'h536;
        15'h0110: data = 12'h46D;
        15'h0111: data = 12'h3A1;
        15'h0112: data = 12'h2EB;
        15'h0113: data = 12'h23F;
        15'h0114: data = 12'h1A5;
        15'h0115: data = 12'h50D;
        15'h0116: data = 12'h0BA;
        15'h0117: data = 12'h056;
        15'h0118: data = 12'h785;
        15'h0119: data = 12'h776;
        15'h011A: data = 12'h777;
        15'h011B: data = 12'h75E;
        15'h011C: data = 12'h785;
        15'h011D: data = 12'h7A6;
        15'h011E: data = 12'h7EA;
        15'h011F: data = 12'h099;
        15'h0120: data = 12'h107;
        15'h0121: data = 12'h176;
        15'h0122: data = 12'h203;
        15'h0123: data = 12'h2A4;
        15'h0124: data = 12'h357;
        15'h0125: data = 12'h41F;
        15'h0126: data = 12'h4F7;
        15'h0127: data = 12'h5DB;
        15'h0128: data = 12'h6CE;
        15'h0129: data = 12'h7C9;
        15'h012A: data = 12'h0FD;
        15'h012B: data = 12'h209;
        15'h012C: data = 12'h313;
        15'h012D: data = 12'h430;
        15'h012E: data = 12'h53D;
        15'h012F: data = 12'h65A;
        15'h0130: data = 12'h782;
        15'h0131: data = 12'h0ED;
        15'h0132: data = 12'h20E;
        15'h0133: data = 12'h332;
        15'h0134: data = 12'h50D;
        15'h0135: data = 12'h55C;
        15'h0136: data = 12'h65E;
        15'h0137: data = 12'h752;
        15'h0138: data = 12'h57C;
        15'h0139: data = 12'h15F;
        15'h013A: data = 12'h230;
        15'h013B: data = 12'h2F2;
        15'h013C: data = 12'h3AF;
        15'h013D: data = 12'h44E;
        15'h013E: data = 12'h4E4;
        15'h013F: data = 12'h559;
        15'h0140: data = 12'h5D1;
        15'h0141: data = 12'h617;
        15'h0142: data = 12'h659;
        15'h0143: data = 12'h687;
        15'h0144: data = 12'h68F;
        15'h0145: data = 12'h684;
        15'h0146: data = 12'h666;
        15'h0147: data = 12'h638;
        15'h0148: data = 12'h5E4;
        15'h0149: data = 12'h59A;
        15'h014A: data = 12'h535;
        15'h014B: data = 12'h4B5;
        15'h014C: data = 12'h41D;
        15'h014D: data = 12'h371;
        15'h014E: data = 12'h2BA;
        15'h014F: data = 12'h1EB;
        15'h0150: data = 12'h10C;
        15'h0151: data = 12'h020;
        15'h0152: data = 12'h6E9;
        15'h0153: data = 12'h50D;
        15'h0154: data = 12'h4E0;
        15'h0155: data = 12'h3D1;
        15'h0156: data = 12'h2B2;
        15'h0157: data = 12'h1A0;
        15'h0158: data = 12'h08C;
        15'h0159: data = 12'h70F;
        15'h015A: data = 12'h5FB;
        15'h015B: data = 12'h4E7;
        15'h015C: data = 12'h3BE;
        15'h015D: data = 12'h2B0;
        15'h015E: data = 12'h18F;
        15'h015F: data = 12'h08A;
        15'h0160: data = 12'h749;
        15'h0161: data = 12'h661;
        15'h0162: data = 12'h573;
        15'h0163: data = 12'h49F;
        15'h0164: data = 12'h3D1;
        15'h0165: data = 12'h31E;
        15'h0166: data = 12'h279;
        15'h0167: data = 12'h1D9;
        15'h0168: data = 12'h14D;
        15'h0169: data = 12'h0E6;
        15'h016A: data = 12'h081;
        15'h016B: data = 12'h034;
        15'h016C: data = 12'h795;
        15'h016D: data = 12'h771;
        15'h016E: data = 12'h753;
        15'h016F: data = 12'h775;
        15'h0170: data = 12'h798;
        15'h0171: data = 12'h7D4;
        15'h0172: data = 12'h50D;
        15'h0173: data = 12'h0E0;
        15'h0174: data = 12'h14E;
        15'h0175: data = 12'h1DB;
        15'h0176: data = 12'h278;
        15'h0177: data = 12'h329;
        15'h0178: data = 12'h3E1;
        15'h0179: data = 12'h4AC;
        15'h017A: data = 12'h580;
        15'h017B: data = 12'h673;
        15'h017C: data = 12'h766;
        15'h017D: data = 12'h0E5;
        15'h017E: data = 12'h1A2;
        15'h017F: data = 12'h2C2;
        15'h0180: data = 12'h3D5;
        15'h0181: data = 12'h4F8;
        15'h0182: data = 12'h609;
        15'h0183: data = 12'h71D;
        15'h0184: data = 12'h46C;
        15'h0185: data = 12'h1A5;
        15'h0186: data = 12'h2C7;
        15'h0187: data = 12'h3E7;
        15'h0188: data = 12'h4FF;
        15'h0189: data = 12'h60F;
        15'h018A: data = 12'h70F;
        15'h018B: data = 12'h802;
        15'h018C: data = 12'h124;
        15'h018D: data = 12'h1F4;
        15'h018E: data = 12'h2B3;
        15'h018F: data = 12'h36C;
        15'h0190: data = 12'h416;
        15'h0191: data = 12'h50D;
        15'h0192: data = 12'h538;
        15'h0193: data = 12'h5A8;
        15'h0194: data = 12'h5F9;
        15'h0195: data = 12'h64C;
        15'h0196: data = 12'h675;
        15'h0197: data = 12'h69A;
        15'h0198: data = 12'h694;
        15'h0199: data = 12'h675;
        15'h019A: data = 12'h64B;
        15'h019B: data = 12'h603;
        15'h019C: data = 12'h5B6;
        15'h019D: data = 12'h54B;
        15'h019E: data = 12'h4D5;
        15'h019F: data = 12'h452;
        15'h01A0: data = 12'h3A8;
        15'h01A1: data = 12'h2FA;
        15'h01A2: data = 12'h234;
        15'h01A3: data = 12'h15A;
        15'h01A4: data = 12'h079;
        15'h01A5: data = 12'h745;
        15'h01A6: data = 12'h645;
        15'h01A7: data = 12'h540;
        15'h01A8: data = 12'h427;
        15'h01A9: data = 12'h318;
        15'h01AA: data = 12'h1FB;
        15'h01AB: data = 12'h0DD;
        15'h01AC: data = 12'h77D;
        15'h01AD: data = 12'h654;
        15'h01AE: data = 12'h53A;
        15'h01AF: data = 12'h427;
        15'h01B0: data = 12'h50D;
        15'h01B1: data = 12'h1F3;
        15'h01B2: data = 12'h0E6;
        15'h01B3: data = 12'h776;
        15'h01B4: data = 12'h6AF;
        15'h01B5: data = 12'h5C3;
        15'h01B6: data = 12'h4E9;
        15'h01B7: data = 12'h414;
        15'h01B8: data = 12'h351;
        15'h01B9: data = 12'h2A2;
        15'h01BA: data = 12'h206;
        15'h01BB: data = 12'h177;
        15'h01BC: data = 12'h104;
        15'h01BD: data = 12'h0A2;
        15'h01BE: data = 12'h049;
        15'h01BF: data = 12'h7A1;
        15'h01C0: data = 12'h77E;
        15'h01C1: data = 12'h75B;
        15'h01C2: data = 12'h774;
        15'h01C3: data = 12'h773;
        15'h01C4: data = 12'h7B2;
        15'h01C5: data = 12'h7F3;
        15'h01C6: data = 12'h0B9;
        15'h01C7: data = 12'h11D;
        15'h01C8: data = 12'h1B0;
        15'h01C9: data = 12'h248;
        15'h01CA: data = 12'h2F5;
        15'h01CB: data = 12'h3AA;
        15'h01CC: data = 12'h471;
        15'h01CD: data = 12'h53D;
        15'h01CE: data = 12'h61B;
        15'h01CF: data = 12'h50D;
        15'h01D0: data = 12'h80C;
        15'h01D1: data = 12'h149;
        15'h01D2: data = 12'h260;
        15'h01D3: data = 12'h37C;
        15'h01D4: data = 12'h495;
        15'h01D5: data = 12'h5AE;
        15'h01D6: data = 12'h6CF;
        15'h01D7: data = 12'h7E1;
        15'h01D8: data = 12'h147;
        15'h01D9: data = 12'h269;
        15'h01DA: data = 12'h37F;
        15'h01DB: data = 12'h499;
        15'h01DC: data = 12'h5A8;
        15'h01DD: data = 12'h6B6;
        15'h01DE: data = 12'h7AA;
        15'h01DF: data = 12'h0D3;
        15'h01E0: data = 12'h1BB;
        15'h01E1: data = 12'h286;
        15'h01E2: data = 12'h33A;
        15'h01E3: data = 12'h3EA;
        15'h01E4: data = 12'h486;
        15'h01E5: data = 12'h509;
        15'h01E6: data = 12'h57A;
        15'h01E7: data = 12'h5E9;
        15'h01E8: data = 12'h637;
        15'h01E9: data = 12'h67E;
        15'h01EA: data = 12'h69A;
        15'h01EB: data = 12'h69A;
        15'h01EC: data = 12'h699;
        15'h01ED: data = 12'h670;
        15'h01EE: data = 12'h50D;
        15'h01EF: data = 12'h5E0;
        15'h01F0: data = 12'h570;
        15'h01F1: data = 12'h504;
        15'h01F2: data = 12'h477;
        15'h01F3: data = 12'h3DC;
        15'h01F4: data = 12'h32C;
        15'h01F5: data = 12'h274;
        15'h01F6: data = 12'h1A2;
        15'h01F7: data = 12'h0C7;
        15'h01F8: data = 12'h782;
        15'h01F9: data = 12'h6AA;
        15'h01FA: data = 12'h5A1;
        15'h01FB: data = 12'h494;
        15'h01FC: data = 12'h374;
        15'h01FD: data = 12'h258;
        15'h01FE: data = 12'h137;
        15'h01FF: data = 12'h02D;
        15'h0200: data = 12'h6B2;
        15'h0201: data = 12'h589;
        15'h0202: data = 12'h47C;
        15'h0203: data = 12'h363;
        15'h0204: data = 12'h24E;
        15'h0205: data = 12'h13C;
        15'h0206: data = 12'h039;
        15'h0207: data = 12'h70B;
        15'h0208: data = 12'h61A;
        15'h0209: data = 12'h533;
        15'h020A: data = 12'h45F;
        15'h020B: data = 12'h391;
        15'h020C: data = 12'h2DB;
        15'h020D: data = 12'h50D;
        15'h020E: data = 12'h19E;
        15'h020F: data = 12'h115;
        15'h0210: data = 12'h0C4;
        15'h0211: data = 12'h063;
        15'h0212: data = 12'h691;
        15'h0213: data = 12'h789;
        15'h0214: data = 12'h77E;
        15'h0215: data = 12'h75D;
        15'h0216: data = 12'h779;
        15'h0217: data = 12'h796;
        15'h0218: data = 12'h7D6;
        15'h0219: data = 12'h091;
        15'h021A: data = 12'h0FC;
        15'h021B: data = 12'h176;
        15'h021C: data = 12'h20D;
        15'h021D: data = 12'h2B7;
        15'h021E: data = 12'h36A;
        15'h021F: data = 12'h432;
        15'h0220: data = 12'h503;
        15'h0221: data = 12'h5E2;
        15'h0222: data = 12'h6C8;
        15'h0223: data = 12'h7C0;
        15'h0224: data = 12'h0ED;
        15'h0225: data = 12'h1F7;
        15'h0226: data = 12'h30A;
        15'h0227: data = 12'h430;
        15'h0228: data = 12'h54A;
        15'h0229: data = 12'h674;
        15'h022A: data = 12'h798;
        15'h022B: data = 12'h0FA;
        15'h022C: data = 12'h50D;
        15'h022D: data = 12'h32F;
        15'h022E: data = 12'h43B;
        15'h022F: data = 12'h54A;
        15'h0230: data = 12'h650;
        15'h0231: data = 12'h74F;
        15'h0232: data = 12'h2D6;
        15'h0233: data = 12'h16F;
        15'h0234: data = 12'h242;
        15'h0235: data = 12'h303;
        15'h0236: data = 12'h3BB;
        15'h0237: data = 12'h457;
        15'h0238: data = 12'h4E5;
        15'h0239: data = 12'h553;
        15'h023A: data = 12'h5C3;
        15'h023B: data = 12'h604;
        15'h023C: data = 12'h648;
        15'h023D: data = 12'h67A;
        15'h023E: data = 12'h690;
        15'h023F: data = 12'h693;
        15'h0240: data = 12'h67A;
        15'h0241: data = 12'h648;
        15'h0242: data = 12'h5F2;
        15'h0243: data = 12'h5A2;
        15'h0244: data = 12'h534;
        15'h0245: data = 12'h4A8;
        15'h0246: data = 12'h40A;
        15'h0247: data = 12'h361;
        15'h0248: data = 12'h2AB;
        15'h0249: data = 12'h1DF;
        15'h024A: data = 12'h10D;
        15'h024B: data = 12'h50D;
        15'h024C: data = 12'h6FA;
        15'h024D: data = 12'h5FE;
        15'h024E: data = 12'h4F4;
        15'h024F: data = 12'h3E0;
        15'h0250: data = 12'h2BF;
        15'h0251: data = 12'h1A4;
        15'h0252: data = 12'h082;
        15'h0253: data = 12'h701;
        15'h0254: data = 12'h5EB;
        15'h0255: data = 12'h4D7;
        15'h0256: data = 12'h3B6;
        15'h0257: data = 12'h2A9;
        15'h0258: data = 12'h196;
        15'h0259: data = 12'h096;
        15'h025A: data = 12'h75B;
        15'h025B: data = 12'h674;
        15'h025C: data = 12'h57E;
        15'h025D: data = 12'h4AB;
        15'h025E: data = 12'h3D4;
        15'h025F: data = 12'h316;
        15'h0260: data = 12'h268;
        15'h0261: data = 12'h1CC;
        15'h0262: data = 12'h140;
        15'h0263: data = 12'h0DA;
        15'h0264: data = 12'h080;
        15'h0265: data = 12'h038;
        15'h0266: data = 12'h7A5;
        15'h0267: data = 12'h789;
        15'h0268: data = 12'h767;
        15'h0269: data = 12'h782;
        15'h026A: data = 12'h50D;
        15'h026B: data = 12'h7D7;
        15'h026C: data = 12'h4E9;
        15'h026D: data = 12'h0D5;
        15'h026E: data = 12'h144;
        15'h026F: data = 12'h1CD;
        15'h0270: data = 12'h272;
        15'h0271: data = 12'h32C;
        15'h0272: data = 12'h3ED;
        15'h0273: data = 12'h4C0;
        15'h0274: data = 12'h596;
        15'h0275: data = 12'h683;
        15'h0276: data = 12'h76D;
        15'h0277: data = 12'h197;
        15'h0278: data = 12'h195;
        15'h0279: data = 12'h2AE;
        15'h027A: data = 12'h3C8;
        15'h027B: data = 12'h4EF;
        15'h027C: data = 12'h60A;
        15'h027D: data = 12'h72C;
        15'h027E: data = 12'h759;
        15'h027F: data = 12'h1B9;
        15'h0280: data = 12'h2D4;
        15'h0281: data = 12'h3EE;
        15'h0282: data = 12'h4F9;
        15'h0283: data = 12'h601;
        15'h0284: data = 12'h6FE;
        15'h0285: data = 12'h7F1;
        15'h0286: data = 12'h115;
        15'h0287: data = 12'h1EB;
        15'h0288: data = 12'h2BC;
        15'h0289: data = 12'h50D;
        15'h028A: data = 12'h425;
        15'h028B: data = 12'h4BC;
        15'h028C: data = 12'h542;
        15'h028D: data = 12'h5A6;
        15'h028E: data = 12'h5EA;
        15'h028F: data = 12'h63C;
        15'h0290: data = 12'h665;
        15'h0291: data = 12'h689;
        15'h0292: data = 12'h68F;
        15'h0293: data = 12'h67B;
        15'h0294: data = 12'h658;
        15'h0295: data = 12'h61B;
        15'h0296: data = 12'h5CF;
        15'h0297: data = 12'h55B;
        15'h0298: data = 12'h4D8;
        15'h0299: data = 12'h44D;
        15'h029A: data = 12'h39F;
        15'h029B: data = 12'h2E9;
        15'h029C: data = 12'h223;
        15'h029D: data = 12'h14A;
        15'h029E: data = 12'h071;
        15'h029F: data = 12'h741;
        15'h02A0: data = 12'h64D;
        15'h02A1: data = 12'h54B;
        15'h02A2: data = 12'h439;
        15'h02A3: data = 12'h329;
        15'h02A4: data = 12'h209;
        15'h02A5: data = 12'h0EC;
        15'h02A6: data = 12'h75F;
        15'h02A7: data = 12'h64C;
        15'h02A8: data = 12'h50D;
        15'h02A9: data = 12'h416;
        15'h02AA: data = 12'h2F8;
        15'h02AB: data = 12'h1E8;
        15'h02AC: data = 12'h0E7;
        15'h02AD: data = 12'h64E;
        15'h02AE: data = 12'h6BE;
        15'h02AF: data = 12'h5D4;
        15'h02B0: data = 12'h4F7;
        15'h02B1: data = 12'h422;
        15'h02B2: data = 12'h35C;
        15'h02B3: data = 12'h2A4;
        15'h02B4: data = 12'h1FD;
        15'h02B5: data = 12'h16F;
        15'h02B6: data = 12'h0F7;
        15'h02B7: data = 12'h099;
        15'h02B8: data = 12'h040;
        15'h02B9: data = 12'h79E;
        15'h02BA: data = 12'h783;
        15'h02BB: data = 12'h764;
        15'h02BC: data = 12'h780;
        15'h02BD: data = 12'h781;
        15'h02BE: data = 12'h7C0;
        15'h02BF: data = 12'h7FB;
        15'h02C0: data = 12'h0BB;
        15'h02C1: data = 12'h113;
        15'h02C2: data = 12'h1A2;
        15'h02C3: data = 12'h236;
        15'h02C4: data = 12'h2E3;
        15'h02C5: data = 12'h3A1;
        15'h02C6: data = 12'h473;
        15'h02C7: data = 12'h50D;
        15'h02C8: data = 12'h635;
        15'h02C9: data = 12'h720;
        15'h02CA: data = 12'h81B;
        15'h02CB: data = 12'h14A;
        15'h02CC: data = 12'h257;
        15'h02CD: data = 12'h36B;
        15'h02CE: data = 12'h482;
        15'h02CF: data = 12'h59F;
        15'h02D0: data = 12'h6CF;
        15'h02D1: data = 12'h7EE;
        15'h02D2: data = 12'h15C;
        15'h02D3: data = 12'h27C;
        15'h02D4: data = 12'h38F;
        15'h02D5: data = 12'h4A2;
        15'h02D6: data = 12'h5A4;
        15'h02D7: data = 12'h6A8;
        15'h02D8: data = 12'h799;
        15'h02D9: data = 12'h0C4;
        15'h02DA: data = 12'h1AA;
        15'h02DB: data = 12'h27C;
        15'h02DC: data = 12'h33D;
        15'h02DD: data = 12'h3F4;
        15'h02DE: data = 12'h497;
        15'h02DF: data = 12'h51A;
        15'h02E0: data = 12'h582;
        15'h02E1: data = 12'h5E7;
        15'h02E2: data = 12'h628;
        15'h02E3: data = 12'h667;
        15'h02E4: data = 12'h683;
        15'h02E5: data = 12'h688;
        15'h02E6: data = 12'h50D;
        15'h02E7: data = 12'h66F;
        15'h02E8: data = 12'h637;
        15'h02E9: data = 12'h5E8;
        15'h02EA: data = 12'h57C;
        15'h02EB: data = 12'h515;
        15'h02EC: data = 12'h482;
        15'h02ED: data = 12'h3DE;
        15'h02EE: data = 12'h32C;
        15'h02EF: data = 12'h269;
        15'h02F0: data = 12'h191;
        15'h02F1: data = 12'h0B3;
        15'h02F2: data = 12'h791;
        15'h02F3: data = 12'h69D;
        15'h02F4: data = 12'h59D;
        15'h02F5: data = 12'h49D;
        15'h02F6: data = 12'h37B;
        15'h02F7: data = 12'h264;
        15'h02F8: data = 12'h143;
        15'h02F9: data = 12'h025;
        15'h02FA: data = 12'h6B5;
        15'h02FB: data = 12'h587;
        15'h02FC: data = 12'h471;
        15'h02FD: data = 12'h354;
        15'h02FE: data = 12'h23D;
        15'h02FF: data = 12'h130;
        15'h0300: data = 12'h030;
        15'h0301: data = 12'h705;
        15'h0302: data = 12'h61E;
        15'h0303: data = 12'h538;
        15'h0304: data = 12'h469;
        15'h0305: data = 12'h50D;
        15'h0306: data = 12'h2E5;
        15'h0307: data = 12'h232;
        15'h0308: data = 12'h19C;
        15'h0309: data = 12'h10D;
        15'h030A: data = 12'h0B7;
        15'h030B: data = 12'h059;
        15'h030C: data = 12'h67F;
        15'h030D: data = 12'h77B;
        15'h030E: data = 12'h77B;
        15'h030F: data = 12'h765;
        15'h0310: data = 12'h787;
        15'h0311: data = 12'h7A5;
        15'h0312: data = 12'h7E5;
        15'h0313: data = 12'h093;
        15'h0314: data = 12'h0F9;
        15'h0315: data = 12'h16A;
        15'h0316: data = 12'h1FF;
        15'h0317: data = 12'h2A4;
        15'h0318: data = 12'h35F;
        15'h0319: data = 12'h42B;
        15'h031A: data = 12'h504;
        15'h031B: data = 12'h5E7;
        15'h031C: data = 12'h6D2;
        15'h031D: data = 12'h7C5;
        15'h031E: data = 12'h0F7;
        15'h031F: data = 12'h1FB;
        15'h0320: data = 12'h306;
        15'h0321: data = 12'h425;
        15'h0322: data = 12'h53C;
        15'h0323: data = 12'h662;
        15'h0324: data = 12'h50D;
        15'h0325: data = 12'h0F4;
        15'h0326: data = 12'h218;
        15'h0327: data = 12'h335;
        15'h0328: data = 12'h44B;
        15'h0329: data = 12'h559;
        15'h032A: data = 12'h657;
        15'h032B: data = 12'h750;
        15'h032C: data = 12'h330;
        15'h032D: data = 12'h15D;
        15'h032E: data = 12'h233;
        15'h032F: data = 12'h2FD;
        15'h0330: data = 12'h3B6;
        15'h0331: data = 12'h45D;
        15'h0332: data = 12'h4ED;
        15'h0333: data = 12'h565;
        15'h0334: data = 12'h5D1;
        15'h0335: data = 12'h60F;
        15'h0336: data = 12'h64C;
        15'h0337: data = 12'h675;
        15'h0338: data = 12'h685;
        15'h0339: data = 12'h688;
        15'h033A: data = 12'h66E;
        15'h033B: data = 12'h645;
        15'h033C: data = 12'h5F5;
        15'h033D: data = 12'h5A8;
        15'h033E: data = 12'h53D;
        15'h033F: data = 12'h4B0;
        15'h0340: data = 12'h413;
        15'h0341: data = 12'h361;
        15'h0342: data = 12'h2A7;
        15'h0343: data = 12'h50D;
        15'h0344: data = 12'h10A;
        15'h0345: data = 12'h03A;
        15'h0346: data = 12'h6EB;
        15'h0347: data = 12'h5F7;
        15'h0348: data = 12'h4EB;
        15'h0349: data = 12'h3DB;
        15'h034A: data = 12'h2C1;
        15'h034B: data = 12'h1A8;
        15'h034C: data = 12'h089;
        15'h034D: data = 12'h712;
        15'h034E: data = 12'h5F3;
        15'h034F: data = 12'h4D8;
        15'h0350: data = 12'h3AC;
        15'h0351: data = 12'h299;
        15'h0352: data = 12'h186;
        15'h0353: data = 12'h085;
        15'h0354: data = 12'h754;
        15'h0355: data = 12'h672;
        15'h0356: data = 12'h582;
        15'h0357: data = 12'h4B1;
        15'h0358: data = 12'h3DC;
        15'h0359: data = 12'h323;
        15'h035A: data = 12'h277;
        15'h035B: data = 12'h1D4;
        15'h035C: data = 12'h143;
        15'h035D: data = 12'h0D7;
        15'h035E: data = 12'h077;
        15'h035F: data = 12'h02C;
        15'h0360: data = 12'h79D;
        15'h0361: data = 12'h77F;
        15'h0362: data = 12'h50D;
        15'h0363: data = 12'h785;
        15'h0364: data = 12'h7A4;
        15'h0365: data = 12'h7DB;
        15'h0366: data = 12'h7B4;
        15'h0367: data = 12'h0DC;
        15'h0368: data = 12'h145;
        15'h0369: data = 12'h1C9;
        15'h036A: data = 12'h267;
        15'h036B: data = 12'h31B;
        15'h036C: data = 12'h3DD;
        15'h036D: data = 12'h4B6;
        15'h036E: data = 12'h597;
        15'h036F: data = 12'h687;
        15'h0370: data = 12'h776;
        15'h0371: data = 12'h0CE;
        15'h0372: data = 12'h1A0;
        15'h0373: data = 12'h2B6;
        15'h0374: data = 12'h3C6;
        15'h0375: data = 12'h4EC;
        15'h0376: data = 12'h600;
        15'h0377: data = 12'h71F;
        15'h0378: data = 12'h53F;
        15'h0379: data = 12'h1BA;
        15'h037A: data = 12'h2D9;
        15'h037B: data = 12'h3F4;
        15'h037C: data = 12'h506;
        15'h037D: data = 12'h609;
        15'h037E: data = 12'h6FE;
        15'h037F: data = 12'h7F0;
        15'h0380: data = 12'h114;
        15'h0381: data = 12'h50D;
        15'h0382: data = 12'h2B8;
        15'h0383: data = 12'h376;
        15'h0384: data = 12'h423;
        15'h0385: data = 12'h4BF;
        15'h0386: data = 12'h541;
        15'h0387: data = 12'h5AE;
        15'h0388: data = 12'h5FA;
        15'h0389: data = 12'h649;
        15'h038A: data = 12'h666;
        15'h038B: data = 12'h68C;
        15'h038C: data = 12'h687;
        15'h038D: data = 12'h66F;
        15'h038E: data = 12'h64E;
        15'h038F: data = 12'h613;
        15'h0390: data = 12'h5CB;
        15'h0391: data = 12'h55D;
        15'h0392: data = 12'h4DE;
        15'h0393: data = 12'h456;
        15'h0394: data = 12'h3A9;
        15'h0395: data = 12'h2EC;
        15'h0396: data = 12'h220;
        15'h0397: data = 12'h14C;
        15'h0398: data = 12'h068;
        15'h0399: data = 12'h73A;
        15'h039A: data = 12'h645;
        15'h039B: data = 12'h543;
        15'h039C: data = 12'h437;
        15'h039D: data = 12'h32A;
        15'h039E: data = 12'h20B;
        15'h039F: data = 12'h0EA;
        15'h03A0: data = 12'h50D;
        15'h03A1: data = 12'h650;
        15'h03A2: data = 12'h52E;
        15'h03A3: data = 12'h417;
        15'h03A4: data = 12'h2F7;
        15'h03A5: data = 12'h1E0;
        15'h03A6: data = 12'h0DB;
        15'h03A7: data = 12'h7AE;
        15'h03A8: data = 12'h6B8;
        15'h03A9: data = 12'h5D0;
        15'h03AA: data = 12'h4F9;
        15'h03AB: data = 12'h423;
        15'h03AC: data = 12'h35E;
        15'h03AD: data = 12'h2AD;
        15'h03AE: data = 12'h204;
        15'h03AF: data = 12'h171;
        15'h03B0: data = 12'h0F9;
        15'h03B1: data = 12'h095;
        15'h03B2: data = 12'h038;
        15'h03B3: data = 12'h795;
        15'h03B4: data = 12'h77D;
        15'h03B5: data = 12'h762;
        15'h03B6: data = 12'h787;
        15'h03B7: data = 12'h785;
        15'h03B8: data = 12'h7C4;
        15'h03B9: data = 12'h801;
        15'h03BA: data = 12'h0BE;
        15'h03BB: data = 12'h117;
        15'h03BC: data = 12'h1A2;
        15'h03BD: data = 12'h239;
        15'h03BE: data = 12'h2E1;
        15'h03BF: data = 12'h50D;
        15'h03C0: data = 12'h473;
        15'h03C1: data = 12'h548;
        15'h03C2: data = 12'h632;
        15'h03C3: data = 12'h71F;
        15'h03C4: data = 12'h81D;
        15'h03C5: data = 12'h153;
        15'h03C6: data = 12'h25D;
        15'h03C7: data = 12'h372;
        15'h03C8: data = 12'h484;
        15'h03C9: data = 12'h59D;
        15'h03CA: data = 12'h6C5;
        15'h03CB: data = 12'h7E1;
        15'h03CC: data = 12'h158;
        15'h03CD: data = 12'h281;
        15'h03CE: data = 12'h396;
        15'h03CF: data = 12'h4AD;
        15'h03D0: data = 12'h5AF;
        15'h03D1: data = 12'h6B3;
        15'h03D2: data = 12'h79E;
        15'h03D3: data = 12'h0CB;
        15'h03D4: data = 12'h1AB;
        15'h03D5: data = 12'h27A;
        15'h03D6: data = 12'h33D;
        15'h03D7: data = 12'h3F5;
        15'h03D8: data = 12'h498;
        15'h03D9: data = 12'h51D;
        15'h03DA: data = 12'h588;
        15'h03DB: data = 12'h5F1;
        15'h03DC: data = 12'h631;
        15'h03DD: data = 12'h66C;
        15'h03DE: data = 12'h50D;
        15'h03DF: data = 12'h688;
        15'h03E0: data = 12'h687;
        15'h03E1: data = 12'h66C;
        15'h03E2: data = 12'h630;
        15'h03E3: data = 12'h5E9;
        15'h03E4: data = 12'h582;
        15'h03E5: data = 12'h510;
        15'h03E6: data = 12'h485;
        15'h03E7: data = 12'h3E4;
        15'h03E8: data = 12'h331;
        15'h03E9: data = 12'h269;
        15'h03EA: data = 12'h190;
        15'h03EB: data = 12'h0B8;
        15'h03EC: data = 12'h790;
        15'h03ED: data = 12'h69F;
        15'h03EE: data = 12'h59C;
        15'h03EF: data = 12'h497;
        15'h03F0: data = 12'h378;
        15'h03F1: data = 12'h264;
        15'h03F2: data = 12'h144;
        15'h03F3: data = 12'h02C;
        15'h03F4: data = 12'h6BB;
        15'h03F5: data = 12'h58B;
        15'h03F6: data = 12'h475;
        15'h03F7: data = 12'h353;
        15'h03F8: data = 12'h23B;
        15'h03F9: data = 12'h128;
        15'h03FA: data = 12'h02C;
        15'h03FB: data = 12'h703;
        15'h03FC: data = 12'h61C;
        15'h03FD: data = 12'h50D;
        15'h03FE: data = 12'h471;
        15'h03FF: data = 12'h3A3;
        15'h0400: data = 12'h2E8;
        15'h0401: data = 12'h238;
        15'h0402: data = 12'h19B;
        15'h0403: data = 12'h10F;
        15'h0404: data = 12'h0B5;
        15'h0405: data = 12'h057;
        15'h0406: data = 12'h79D;
        15'h0407: data = 12'h77B;
        15'h0408: data = 12'h776;
        15'h0409: data = 12'h760;
        15'h040A: data = 12'h782;
        15'h040B: data = 12'h7A5;
        15'h040C: data = 12'h7EC;
        15'h040D: data = 12'h09C;
        15'h040E: data = 12'h0FF;
        15'h040F: data = 12'h170;
        15'h0410: data = 12'h204;
        15'h0411: data = 12'h2A8;
        15'h0412: data = 12'h35B;
        15'h0413: data = 12'h42B;
        15'h0414: data = 12'h502;
        15'h0415: data = 12'h5E9;
        15'h0416: data = 12'h6D2;
        15'h0417: data = 12'h7C9;
        15'h0418: data = 12'h0FD;
        15'h0419: data = 12'h204;
        15'h041A: data = 12'h30E;
        15'h041B: data = 12'h42A;
        15'h041C: data = 12'h50D;
        15'h041D: data = 12'h665;
        15'h041E: data = 12'h787;
        15'h041F: data = 12'h0F8;
        15'h0420: data = 12'h217;
        15'h0421: data = 12'h341;
        15'h0422: data = 12'h44C;
        15'h0423: data = 12'h55D;
        15'h0424: data = 12'h65C;
        15'h0425: data = 12'h750;
        15'h0426: data = 12'h339;
        15'h0427: data = 12'h15F;
        15'h0428: data = 12'h233;
        15'h0429: data = 12'h303;
        15'h042A: data = 12'h3BC;
        15'h042B: data = 12'h460;
        15'h042C: data = 12'h4EF;
        15'h042D: data = 12'h562;
        15'h042E: data = 12'h5D0;
        15'h042F: data = 12'h615;
        15'h0430: data = 12'h64E;
        15'h0431: data = 12'h678;
        15'h0432: data = 12'h68B;
        15'h0433: data = 12'h68E;
        15'h0434: data = 12'h669;
        15'h0435: data = 12'h643;
        15'h0436: data = 12'h5F8;
        15'h0437: data = 12'h5A6;
        15'h0438: data = 12'h542;
        15'h0439: data = 12'h4B4;
        15'h043A: data = 12'h417;
        15'h043B: data = 12'h50D;
        15'h043C: data = 12'h2AB;
        15'h043D: data = 12'h1DA;
        15'h043E: data = 12'h102;
        15'h043F: data = 12'h036;
        15'h0440: data = 12'h6EB;
        15'h0441: data = 12'h5F7;
        15'h0442: data = 12'h4EC;
        15'h0443: data = 12'h3E3;
        15'h0444: data = 12'h2C1;
        15'h0445: data = 12'h1A9;
        15'h0446: data = 12'h08C;
        15'h0447: data = 12'h70A;
        15'h0448: data = 12'h5F7;
        15'h0449: data = 12'h4D5;
        15'h044A: data = 12'h3AE;
        15'h044B: data = 12'h29D;
        15'h044C: data = 12'h184;
        15'h044D: data = 12'h08A;
        15'h044E: data = 12'h751;
        15'h044F: data = 12'h66D;
        15'h0450: data = 12'h57F;
        15'h0451: data = 12'h4B1;
        15'h0452: data = 12'h3DC;
        15'h0453: data = 12'h320;
        15'h0454: data = 12'h276;
        15'h0455: data = 12'h1D3;
        15'h0456: data = 12'h13E;
        15'h0457: data = 12'h0D9;
        15'h0458: data = 12'h074;
        15'h0459: data = 12'h02B;
        15'h045A: data = 12'h50D;
        15'h045B: data = 12'h77E;
        15'h045C: data = 12'h764;
        15'h045D: data = 12'h786;
        15'h045E: data = 12'h7A9;
        15'h045F: data = 12'h7E1;
        15'h0460: data = 12'h752;
        15'h0461: data = 12'h0DD;
        15'h0462: data = 12'h140;
        15'h0463: data = 12'h1CE;
        15'h0464: data = 12'h271;
        15'h0465: data = 12'h323;
        15'h0466: data = 12'h3E3;
        15'h0467: data = 12'h4B7;
        15'h0468: data = 12'h595;
        15'h0469: data = 12'h686;
        15'h046A: data = 12'h772;
        15'h046B: data = 12'h0D4;
        15'h046C: data = 12'h1A6;
        15'h046D: data = 12'h2BC;
        15'h046E: data = 12'h3C9;
        15'h046F: data = 12'h4EB;
        15'h0470: data = 12'h601;
        15'h0471: data = 12'h71D;
        15'h0472: data = 12'h478;
        15'h0473: data = 12'h1B9;
        15'h0474: data = 12'h2DC;
        15'h0475: data = 12'h3FB;
        15'h0476: data = 12'h509;
        15'h0477: data = 12'h60A;
        15'h0478: data = 12'h701;
        15'h0479: data = 12'h50D;
        15'h047A: data = 12'h115;
        15'h047B: data = 12'h1EA;
        15'h047C: data = 12'h2BC;
        15'h047D: data = 12'h377;
        15'h047E: data = 12'h427;
        15'h047F: data = 12'h4C0;
        15'h0480: data = 12'h546;
        15'h0481: data = 12'h5AF;
        15'h0482: data = 12'h5F3;
        15'h0483: data = 12'h646;
        15'h0484: data = 12'h66D;
        15'h0485: data = 12'h684;
        15'h0486: data = 12'h688;
        15'h0487: data = 12'h674;
        15'h0488: data = 12'h653;
        15'h0489: data = 12'h616;
        15'h048A: data = 12'h5CA;
        15'h048B: data = 12'h55E;
        15'h048C: data = 12'h4E1;
        15'h048D: data = 12'h45A;
        15'h048E: data = 12'h3A7;
        15'h048F: data = 12'h2EA;
        15'h0490: data = 12'h221;
        15'h0491: data = 12'h14B;
        15'h0492: data = 12'h06C;
        15'h0493: data = 12'h734;
        15'h0494: data = 12'h644;
        15'h0495: data = 12'h547;
        15'h0496: data = 12'h438;
        15'h0497: data = 12'h329;
        15'h0498: data = 12'h50D;
        15'h0499: data = 12'h0EE;
        15'h049A: data = 12'h768;
        15'h049B: data = 12'h651;
        15'h049C: data = 12'h52D;
        15'h049D: data = 12'h413;
        15'h049E: data = 12'h2F5;
        15'h049F: data = 12'h1E0;
        15'h04A0: data = 12'h0DC;
        15'h04A1: data = 12'h7AE;
        15'h04A2: data = 12'h6B5;
        15'h04A3: data = 12'h5D2;
        15'h04A4: data = 12'h4F9;
        15'h04A5: data = 12'h420;
        15'h04A6: data = 12'h35C;
        15'h04A7: data = 12'h2A9;
        15'h04A8: data = 12'h206;
        15'h04A9: data = 12'h176;
        15'h04AA: data = 12'h0FB;
        15'h04AB: data = 12'h094;
        15'h04AC: data = 12'h03A;
        15'h04AD: data = 12'h796;
        15'h04AE: data = 12'h779;
        15'h04AF: data = 12'h75A;
        15'h04B0: data = 12'h77D;
        15'h04B1: data = 12'h785;
        15'h04B2: data = 12'h7C2;
        15'h04B3: data = 12'h801;
        15'h04B4: data = 12'h0C3;
        15'h04B5: data = 12'h11D;
        15'h04B6: data = 12'h1A3;
        15'h04B7: data = 12'h50D;
        15'h04B8: data = 12'h2E1;
        15'h04B9: data = 12'h39A;
        15'h04BA: data = 12'h46C;
        15'h04BB: data = 12'h547;
        15'h04BC: data = 12'h634;
        15'h04BD: data = 12'h720;
        15'h04BE: data = 12'h81E;
        15'h04BF: data = 12'h151;
        15'h04C0: data = 12'h25E;
        15'h04C1: data = 12'h374;
        15'h04C2: data = 12'h486;
        15'h04C3: data = 12'h59C;
        15'h04C4: data = 12'h6C7;
        15'h04C5: data = 12'h7E1;
        15'h04C6: data = 12'h155;
        15'h04C7: data = 12'h27A;
        15'h04C8: data = 12'h393;
        15'h04C9: data = 12'h4AE;
        15'h04CA: data = 12'h5B5;
        15'h04CB: data = 12'h6BD;
        15'h04CC: data = 12'h7A7;
        15'h04CD: data = 12'h0D1;
        15'h04CE: data = 12'h1AE;
        15'h04CF: data = 12'h277;
        15'h04D0: data = 12'h332;
        15'h04D1: data = 12'h3EB;
        15'h04D2: data = 12'h492;
        15'h04D3: data = 12'h51E;
        15'h04D4: data = 12'h58D;
        15'h04D5: data = 12'h5F6;
        15'h04D6: data = 12'h50D;
        15'h04D7: data = 12'h670;
        15'h04D8: data = 12'h68A;
        15'h04D9: data = 12'h687;
        15'h04DA: data = 12'h684;
        15'h04DB: data = 12'h668;
        15'h04DC: data = 12'h62F;
        15'h04DD: data = 12'h5E1;
        15'h04DE: data = 12'h579;
        15'h04DF: data = 12'h512;
        15'h04E0: data = 12'h482;
        15'h04E1: data = 12'h3E5;
        15'h04E2: data = 12'h334;
        15'h04E3: data = 12'h26F;
        15'h04E4: data = 12'h199;
        15'h04E5: data = 12'h0BB;
        15'h04E6: data = 12'h78C;
        15'h04E7: data = 12'h697;
        15'h04E8: data = 12'h592;
        15'h04E9: data = 12'h48D;
        15'h04EA: data = 12'h374;
        15'h04EB: data = 12'h266;
        15'h04EC: data = 12'h14A;
        15'h04ED: data = 12'h02D;
        15'h04EE: data = 12'h6C1;
        15'h04EF: data = 12'h598;
        15'h04F0: data = 12'h480;
        15'h04F1: data = 12'h35B;
        15'h04F2: data = 12'h241;
        15'h04F3: data = 12'h127;
        15'h04F4: data = 12'h029;
        15'h04F5: data = 12'h50D;
        15'h04F6: data = 12'h612;
        15'h04F7: data = 12'h537;
        15'h04F8: data = 12'h468;
        15'h04F9: data = 12'h39C;
        15'h04FA: data = 12'h2E6;
        15'h04FB: data = 12'h23C;
        15'h04FC: data = 12'h1AA;
        15'h04FD: data = 12'h116;
        15'h04FE: data = 12'h0BE;
        15'h04FF: data = 12'h05B;
        15'h0500: data = 12'h7A2;
        15'h0501: data = 12'h772;
        15'h0502: data = 12'h76E;
        15'h0503: data = 12'h75A;
        15'h0504: data = 12'h780;
        15'h0505: data = 12'h7A4;
        15'h0506: data = 12'h7EA;
        15'h0507: data = 12'h09A;
        15'h0508: data = 12'h103;
        15'h0509: data = 12'h177;
        15'h050A: data = 12'h206;
        15'h050B: data = 12'h2A6;
        15'h050C: data = 12'h35B;
        15'h050D: data = 12'h424;
        15'h050E: data = 12'h4F4;
        15'h050F: data = 12'h5DB;
        15'h0510: data = 12'h6CE;
        15'h0511: data = 12'h7CB;
        15'h0512: data = 12'h100;
        15'h0513: data = 12'h207;
        15'h0514: data = 12'h50D;
        15'h0515: data = 12'h431;
        15'h0516: data = 12'h53E;
        15'h0517: data = 12'h663;
        15'h0518: data = 12'h784;
        15'h0519: data = 12'h0F2;
        15'h051A: data = 12'h20C;
        15'h051B: data = 12'h338;
        15'h051C: data = 12'h44E;
        15'h051D: data = 12'h559;
        15'h051E: data = 12'h663;
        15'h051F: data = 12'h75E;
        15'h0520: data = 12'h547;
        15'h0521: data = 12'h167;
        15'h0522: data = 12'h232;
        15'h0523: data = 12'h2F4;
        15'h0524: data = 12'h3AC;
        15'h0525: data = 12'h450;
        15'h0526: data = 12'h4E5;
        15'h0527: data = 12'h55B;
        15'h0528: data = 12'h5D4;
        15'h0529: data = 12'h618;
        15'h052A: data = 12'h659;
        15'h052B: data = 12'h682;
        15'h052C: data = 12'h68C;
        15'h052D: data = 12'h688;
        15'h052E: data = 12'h661;
        15'h052F: data = 12'h62F;
        15'h0530: data = 12'h5E3;
        15'h0531: data = 12'h593;
        15'h0532: data = 12'h532;
        15'h0533: data = 12'h50D;
        15'h0534: data = 12'h41B;
        15'h0535: data = 12'h370;
        15'h0536: data = 12'h2B6;
        15'h0537: data = 12'h1E9;
        15'h0538: data = 12'h108;
        15'h0539: data = 12'h01C;
        15'h053A: data = 12'h6E4;
        15'h053B: data = 12'h5E6;
        15'h053C: data = 12'h4DC;
        15'h053D: data = 12'h3C9;
        15'h053E: data = 12'h2AF;
        15'h053F: data = 12'h19F;
        15'h0540: data = 12'h088;
        15'h0541: data = 12'h70E;
        15'h0542: data = 12'h600;
        15'h0543: data = 12'h4E8;
        15'h0544: data = 12'h3C1;
        15'h0545: data = 12'h2A8;
        15'h0546: data = 12'h186;
        15'h0547: data = 12'h084;
        15'h0548: data = 12'h748;
        15'h0549: data = 12'h65D;
        15'h054A: data = 12'h570;
        15'h054B: data = 12'h49F;
        15'h054C: data = 12'h3D3;
        15'h054D: data = 12'h31C;
        15'h054E: data = 12'h277;
        15'h054F: data = 12'h1DE;
        15'h0550: data = 12'h14D;
        15'h0551: data = 12'h0E6;
        15'h0552: data = 12'h50D;
        15'h0553: data = 12'h038;
        15'h0554: data = 12'h79B;
        15'h0555: data = 12'h775;
        15'h0556: data = 12'h74F;
        15'h0557: data = 12'h772;
        15'h0558: data = 12'h797;
        15'h0559: data = 12'h7D6;
        15'h055A: data = 12'h81F;
        15'h055B: data = 12'h0E4;
        15'h055C: data = 12'h156;
        15'h055D: data = 12'h1DD;
        15'h055E: data = 12'h27B;
        15'h055F: data = 12'h326;
        15'h0560: data = 12'h3DE;
        15'h0561: data = 12'h4A6;
        15'h0562: data = 12'h57F;
        15'h0563: data = 12'h674;
        15'h0564: data = 12'h767;
        15'h0565: data = 12'h0FC;
        15'h0566: data = 12'h1A2;
        15'h0567: data = 12'h2C6;
        15'h0568: data = 12'h3D5;
        15'h0569: data = 12'h4FA;
        15'h056A: data = 12'h60A;
        15'h056B: data = 12'h71B;
        15'h056C: data = 12'h479;
        15'h056D: data = 12'h1A9;
        15'h056E: data = 12'h2C9;
        15'h056F: data = 12'h3EA;
        15'h0570: data = 12'h502;
        15'h0571: data = 12'h50D;
        15'h0572: data = 12'h70D;
        15'h0573: data = 12'h7FD;
        15'h0574: data = 12'h120;
        15'h0575: data = 12'h1F3;
        15'h0576: data = 12'h2B6;
        15'h0577: data = 12'h36C;
        15'h0578: data = 12'h411;
        15'h0579: data = 12'h4AB;
        15'h057A: data = 12'h533;
        15'h057B: data = 12'h5A3;
        15'h057C: data = 12'h5FA;
        15'h057D: data = 12'h64F;
        15'h057E: data = 12'h676;
        15'h057F: data = 12'h698;
        15'h0580: data = 12'h68F;
        15'h0581: data = 12'h670;
        15'h0582: data = 12'h648;
        15'h0583: data = 12'h603;
        15'h0584: data = 12'h5B6;
        15'h0585: data = 12'h54D;
        15'h0586: data = 12'h4D2;
        15'h0587: data = 12'h44F;
        15'h0588: data = 12'h3A9;
        15'h0589: data = 12'h2F6;
        15'h058A: data = 12'h230;
        15'h058B: data = 12'h15B;
        15'h058C: data = 12'h07A;
        15'h058D: data = 12'h73E;
        15'h058E: data = 12'h642;
        15'h058F: data = 12'h53D;
        15'h0590: data = 12'h50D;
        15'h0591: data = 12'h312;
        15'h0592: data = 12'h1F9;
        15'h0593: data = 12'h0DF;
        15'h0594: data = 12'h779;
        15'h0595: data = 12'h655;
        15'h0596: data = 12'h534;
        15'h0597: data = 12'h429;
        15'h0598: data = 12'h301;
        15'h0599: data = 12'h1EE;
        15'h059A: data = 12'h0E6;
        15'h059B: data = 12'h785;
        15'h059C: data = 12'h6AF;
        15'h059D: data = 12'h5BB;
        15'h059E: data = 12'h4E0;
        15'h059F: data = 12'h40C;
        15'h05A0: data = 12'h349;
        15'h05A1: data = 12'h29E;
        15'h05A2: data = 12'h1FE;
        15'h05A3: data = 12'h176;
        15'h05A4: data = 12'h105;
        15'h05A5: data = 12'h0A2;
        15'h05A6: data = 12'h043;
        15'h05A7: data = 12'h79E;
        15'h05A8: data = 12'h77C;
        15'h05A9: data = 12'h759;
        15'h05AA: data = 12'h76F;
        15'h05AB: data = 12'h772;
        15'h05AC: data = 12'h7AD;
        15'h05AD: data = 12'h7F1;
        15'h05AE: data = 12'h0BA;
        15'h05AF: data = 12'h50D;
        15'h05B0: data = 12'h1B5;
        15'h05B1: data = 12'h247;
        15'h05B2: data = 12'h2F5;
        15'h05B3: data = 12'h3A7;
        15'h05B4: data = 12'h472;
        15'h05B5: data = 12'h541;
        15'h05B6: data = 12'h61C;
        15'h05B7: data = 12'h708;
        15'h05B8: data = 12'h80E;
        15'h05B9: data = 12'h144;
        15'h05BA: data = 12'h25C;
        15'h05BB: data = 12'h37A;
        15'h05BC: data = 12'h499;
        15'h05BD: data = 12'h5AF;
        15'h05BE: data = 12'h6D2;
        15'h05BF: data = 12'h7E9;
        15'h05C0: data = 12'h14F;
        15'h05C1: data = 12'h272;
        15'h05C2: data = 12'h383;
        15'h05C3: data = 12'h49E;
        15'h05C4: data = 12'h5A3;
        15'h05C5: data = 12'h6B3;
        15'h05C6: data = 12'h7AA;
        15'h05C7: data = 12'h0DD;
        15'h05C8: data = 12'h1B8;
        15'h05C9: data = 12'h284;
        15'h05CA: data = 12'h33C;
        15'h05CB: data = 12'h3F0;
        15'h05CC: data = 12'h484;
        15'h05CD: data = 12'h50C;
        15'h05CE: data = 12'h50D;
        15'h05CF: data = 12'h5E1;
        15'h05D0: data = 12'h628;
        15'h05D1: data = 12'h66F;
        15'h05D2: data = 12'h693;
        15'h05D3: data = 12'h696;
        15'h05D4: data = 12'h695;
        15'h05D5: data = 12'h66E;
        15'h05D6: data = 12'h62E;
        15'h05D7: data = 12'h5DB;
        15'h05D8: data = 12'h567;
        15'h05D9: data = 12'h4FC;
        15'h05DA: data = 12'h470;
        15'h05DB: data = 12'h3D8;
        15'h05DC: data = 12'h32C;
        15'h05DD: data = 12'h26F;
        15'h05DE: data = 12'h19E;
        15'h05DF: data = 12'h0C5;
        15'h05E0: data = 12'h795;
        15'h05E1: data = 12'h6A6;
        15'h05E2: data = 12'h59A;
        15'h05E3: data = 12'h48D;
        15'h05E4: data = 12'h36D;
        15'h05E5: data = 12'h251;
        15'h05E6: data = 12'h135;
        15'h05E7: data = 12'h01D;
        15'h05E8: data = 12'h6AC;
        15'h05E9: data = 12'h588;
        15'h05EA: data = 12'h477;
        15'h05EB: data = 12'h35D;
        15'h05EC: data = 12'h249;
        15'h05ED: data = 12'h50D;
        15'h05EE: data = 12'h039;
        15'h05EF: data = 12'h70B;
        15'h05F0: data = 12'h618;
        15'h05F1: data = 12'h533;
        15'h05F2: data = 12'h45D;
        15'h05F3: data = 12'h38D;
        15'h05F4: data = 12'h2D3;
        15'h05F5: data = 12'h22C;
        15'h05F6: data = 12'h198;
        15'h05F7: data = 12'h116;
        15'h05F8: data = 12'h0C0;
        15'h05F9: data = 12'h067;
        15'h05FA: data = 12'h6C0;
        15'h05FB: data = 12'h783;
        15'h05FC: data = 12'h77C;
        15'h05FD: data = 12'h75C;
        15'h05FE: data = 12'h777;
        15'h05FF: data = 12'h796;
        15'h0600: data = 12'h7DA;
        15'h0601: data = 12'h098;
        15'h0602: data = 12'h0FD;
        15'h0603: data = 12'h177;
        15'h0604: data = 12'h20A;
        15'h0605: data = 12'h2B3;
        15'h0606: data = 12'h367;
        15'h0607: data = 12'h431;
        15'h0608: data = 12'h504;
        15'h0609: data = 12'h5E4;
        15'h060A: data = 12'h6C4;
        15'h060B: data = 12'h7BC;
        15'h060C: data = 12'h50D;
        15'h060D: data = 12'h1F7;
        15'h060E: data = 12'h308;
        15'h060F: data = 12'h431;
        15'h0610: data = 12'h54A;
        15'h0611: data = 12'h670;
        15'h0612: data = 12'h791;
        15'h0613: data = 12'h0F6;
        15'h0614: data = 12'h212;
        15'h0615: data = 12'h333;
        15'h0616: data = 12'h441;
        15'h0617: data = 12'h54D;
        15'h0618: data = 12'h651;
        15'h0619: data = 12'h752;
        15'h061A: data = 12'h3F7;
        15'h061B: data = 12'h16A;
        15'h061C: data = 12'h242;
        15'h061D: data = 12'h301;
        15'h061E: data = 12'h3B8;
        15'h061F: data = 12'h456;
        15'h0620: data = 12'h4E4;
        15'h0621: data = 12'h551;
        15'h0622: data = 12'h5C0;
        15'h0623: data = 12'h603;
        15'h0624: data = 12'h64A;
        15'h0625: data = 12'h67B;
        15'h0626: data = 12'h691;
        15'h0627: data = 12'h695;
        15'h0628: data = 12'h672;
        15'h0629: data = 12'h644;
        15'h062A: data = 12'h5F1;
        15'h062B: data = 12'h50D;
        15'h062C: data = 12'h52D;
        15'h062D: data = 12'h49F;
        15'h062E: data = 12'h40B;
        15'h062F: data = 12'h35F;
        15'h0630: data = 12'h2AA;
        15'h0631: data = 12'h1DE;
        15'h0632: data = 12'h10C;
        15'h0633: data = 12'h080;
        15'h0634: data = 12'h6F0;
        15'h0635: data = 12'h5F5;
        15'h0636: data = 12'h4EB;
        15'h0637: data = 12'h3D7;
        15'h0638: data = 12'h2BB;
        15'h0639: data = 12'h19A;
        15'h063A: data = 12'h077;
        15'h063B: data = 12'h704;
        15'h063C: data = 12'h5ED;
        15'h063D: data = 12'h4D4;
        15'h063E: data = 12'h3B0;
        15'h063F: data = 12'h2A2;
        15'h0640: data = 12'h18F;
        15'h0641: data = 12'h092;
        15'h0642: data = 12'h757;
        15'h0643: data = 12'h670;
        15'h0644: data = 12'h57E;
        15'h0645: data = 12'h4A3;
        15'h0646: data = 12'h3CF;
        15'h0647: data = 12'h310;
        15'h0648: data = 12'h267;
        15'h0649: data = 12'h1C5;
        15'h064A: data = 12'h50D;
        15'h064B: data = 12'h0D4;
        15'h064C: data = 12'h07B;
        15'h064D: data = 12'h037;
        15'h064E: data = 12'h7A4;
        15'h064F: data = 12'h786;
        15'h0650: data = 12'h762;
        15'h0651: data = 12'h780;
        15'h0652: data = 12'h79D;
        15'h0653: data = 12'h7D0;
        15'h0654: data = 12'h558;
        15'h0655: data = 12'h0D3;
        15'h0656: data = 12'h143;
        15'h0657: data = 12'h1D1;
        15'h0658: data = 12'h27B;
        15'h0659: data = 12'h330;
        15'h065A: data = 12'h3EC;
        15'h065B: data = 12'h4C1;
        15'h065C: data = 12'h590;
        15'h065D: data = 12'h683;
        15'h065E: data = 12'h76F;
        15'h065F: data = 12'h1C3;
        15'h0660: data = 12'h195;
        15'h0661: data = 12'h2B4;
        15'h0662: data = 12'h3CB;
        15'h0663: data = 12'h4F2;
        15'h0664: data = 12'h60C;
        15'h0665: data = 12'h72B;
        15'h0666: data = 12'h74E;
        15'h0667: data = 12'h1BD;
        15'h0668: data = 12'h2D8;
        15'h0669: data = 12'h50D;
        15'h066A: data = 12'h4FB;
        15'h066B: data = 12'h5FB;
        15'h066C: data = 12'h6FA;
        15'h066D: data = 12'h7EE;
        15'h066E: data = 12'h119;
        15'h066F: data = 12'h1F2;
        15'h0670: data = 12'h2C5;
        15'h0671: data = 12'h381;
        15'h0672: data = 12'h427;
        15'h0673: data = 12'h4BC;
        15'h0674: data = 12'h53D;
        15'h0675: data = 12'h5A0;
        15'h0676: data = 12'h5EA;
        15'h0677: data = 12'h63F;
        15'h0678: data = 12'h66A;
        15'h0679: data = 12'h68F;
        15'h067A: data = 12'h690;
        15'h067B: data = 12'h676;
        15'h067C: data = 12'h655;
        15'h067D: data = 12'h616;
        15'h067E: data = 12'h5C6;
        15'h067F: data = 12'h557;
        15'h0680: data = 12'h4D9;
        15'h0681: data = 12'h448;
        15'h0682: data = 12'h39B;
        15'h0683: data = 12'h2E6;
        15'h0684: data = 12'h21C;
        15'h0685: data = 12'h146;
        15'h0686: data = 12'h06B;
        15'h0687: data = 12'h742;
        15'h0688: data = 12'h50D;
        15'h0689: data = 12'h54E;
        15'h068A: data = 12'h436;
        15'h068B: data = 12'h32A;
        15'h068C: data = 12'h206;
        15'h068D: data = 12'h0E2;
        15'h068E: data = 12'h76C;
        15'h068F: data = 12'h646;
        15'h0690: data = 12'h525;
        15'h0691: data = 12'h40F;
        15'h0692: data = 12'h2FB;
        15'h0693: data = 12'h1E1;
        15'h0694: data = 12'h0E0;
        15'h0695: data = 12'h7B6;
        15'h0696: data = 12'h6B8;
        15'h0697: data = 12'h5D4;
        15'h0698: data = 12'h4FB;
        15'h0699: data = 12'h420;
        15'h069A: data = 12'h35B;
        15'h069B: data = 12'h2A3;
        15'h069C: data = 12'h1F9;
        15'h069D: data = 12'h16A;
        15'h069E: data = 12'h0F7;
        15'h069F: data = 12'h097;
        15'h06A0: data = 12'h03D;
        15'h06A1: data = 12'h79C;
        15'h06A2: data = 12'h783;
        15'h06A3: data = 12'h766;
        15'h06A4: data = 12'h783;
        15'h06A5: data = 12'h787;
        15'h06A6: data = 12'h7C1;
        15'h06A7: data = 12'h50D;
        15'h06A8: data = 12'h0BB;
        15'h06A9: data = 12'h116;
        15'h06AA: data = 12'h1A1;
        15'h06AB: data = 12'h238;
        15'h06AC: data = 12'h2E3;
        15'h06AD: data = 12'h3A2;
        15'h06AE: data = 12'h477;
        15'h06AF: data = 12'h551;
        15'h06B0: data = 12'h639;
        15'h06B1: data = 12'h722;
        15'h06B2: data = 12'h820;
        15'h06B3: data = 12'h14A;
        15'h06B4: data = 12'h256;
        15'h06B5: data = 12'h36D;
        15'h06B6: data = 12'h48B;
        15'h06B7: data = 12'h5A0;
        15'h06B8: data = 12'h6D0;
        15'h06B9: data = 12'h7ED;
        15'h06BA: data = 12'h15E;
        15'h06BB: data = 12'h280;
        15'h06BC: data = 12'h396;
        15'h06BD: data = 12'h4AE;
        15'h06BE: data = 12'h5A8;
        15'h06BF: data = 12'h6B4;
        15'h06C0: data = 12'h7A0;
        15'h06C1: data = 12'h0D0;
        15'h06C2: data = 12'h1A7;
        15'h06C3: data = 12'h281;
        15'h06C4: data = 12'h342;
        15'h06C5: data = 12'h3F8;
        15'h06C6: data = 12'h50D;
        15'h06C7: data = 12'h51E;
        15'h06C8: data = 12'h58A;
        15'h06C9: data = 12'h5EA;
        15'h06CA: data = 12'h629;
        15'h06CB: data = 12'h669;
        15'h06CC: data = 12'h68C;
        15'h06CD: data = 12'h689;
        15'h06CE: data = 12'h689;
        15'h06CF: data = 12'h66D;
        15'h06D0: data = 12'h634;
        15'h06D1: data = 12'h5E5;
        15'h06D2: data = 12'h57B;
        15'h06D3: data = 12'h50D;
        15'h06D4: data = 12'h482;
        15'h06D5: data = 12'h3E1;
        15'h06D6: data = 12'h32D;
        15'h06D7: data = 12'h268;
        15'h06D8: data = 12'h194;
        15'h06D9: data = 12'h0B9;
        15'h06DA: data = 12'h795;
        15'h06DB: data = 12'h69D;
        15'h06DC: data = 12'h59B;
        15'h06DD: data = 12'h49A;
        15'h06DE: data = 12'h381;
        15'h06DF: data = 12'h26A;
        15'h06E0: data = 12'h146;
        15'h06E1: data = 12'h027;
        15'h06E2: data = 12'h6B4;
        15'h06E3: data = 12'h589;
        15'h06E4: data = 12'h474;
        15'h06E5: data = 12'h50D;
        15'h06E6: data = 12'h23A;
        15'h06E7: data = 12'h12B;
        15'h06E8: data = 12'h02D;
        15'h06E9: data = 12'h702;
        15'h06EA: data = 12'h61A;
        15'h06EB: data = 12'h53B;
        15'h06EC: data = 12'h46A;
        15'h06ED: data = 12'h39B;
        15'h06EE: data = 12'h2E1;
        15'h06EF: data = 12'h237;
        15'h06F0: data = 12'h19A;
        15'h06F1: data = 12'h10D;
        15'h06F2: data = 12'h0B7;
        15'h06F3: data = 12'h059;
        15'h06F4: data = 12'h7BC;
        15'h06F5: data = 12'h778;
        15'h06F6: data = 12'h777;
        15'h06F7: data = 12'h762;
        15'h06F8: data = 12'h786;
        15'h06F9: data = 12'h7A8;
        15'h06FA: data = 12'h7E7;
        15'h06FB: data = 12'h099;
        15'h06FC: data = 12'h0FF;
        15'h06FD: data = 12'h16E;
        15'h06FE: data = 12'h1FD;
        15'h06FF: data = 12'h2A4;
        15'h0700: data = 12'h35C;
        15'h0701: data = 12'h42E;
        15'h0702: data = 12'h508;
        15'h0703: data = 12'h5EC;
        15'h0704: data = 12'h50D;
        15'h0705: data = 12'h7CC;
        15'h0706: data = 12'h0FC;
        15'h0707: data = 12'h1FD;
        15'h0708: data = 12'h307;
        15'h0709: data = 12'h428;
        15'h070A: data = 12'h53A;
        15'h070B: data = 12'h665;
        15'h070C: data = 12'h794;
        15'h070D: data = 12'h101;
        15'h070E: data = 12'h219;
        15'h070F: data = 12'h33C;
        15'h0710: data = 12'h44D;
        15'h0711: data = 12'h559;
        15'h0712: data = 12'h65D;
        15'h0713: data = 12'h752;
        15'h0714: data = 12'h2D5;
        15'h0715: data = 12'h167;
        15'h0716: data = 12'h237;
        15'h0717: data = 12'h2FE;
        15'h0718: data = 12'h3BC;
        15'h0719: data = 12'h45E;
        15'h071A: data = 12'h4F2;
        15'h071B: data = 12'h564;
        15'h071C: data = 12'h5D3;
        15'h071D: data = 12'h60E;
        15'h071E: data = 12'h648;
        15'h071F: data = 12'h676;
        15'h0720: data = 12'h687;
        15'h0721: data = 12'h684;
        15'h0722: data = 12'h66A;
        15'h0723: data = 12'h50D;
        15'h0724: data = 12'h5F5;
        15'h0725: data = 12'h5A3;
        15'h0726: data = 12'h53A;
        15'h0727: data = 12'h4B2;
        15'h0728: data = 12'h416;
        15'h0729: data = 12'h361;
        15'h072A: data = 12'h2A9;
        15'h072B: data = 12'h1D6;
        15'h072C: data = 12'h104;
        15'h072D: data = 12'h037;
        15'h072E: data = 12'h6ED;
        15'h072F: data = 12'h5F3;
        15'h0730: data = 12'h4EA;
        15'h0731: data = 12'h3D8;
        15'h0732: data = 12'h2C1;
        15'h0733: data = 12'h1A6;
        15'h0734: data = 12'h087;
        15'h0735: data = 12'h70E;
        15'h0736: data = 12'h5F5;
        15'h0737: data = 12'h4DA;
        15'h0738: data = 12'h3AD;
        15'h0739: data = 12'h298;
        15'h073A: data = 12'h180;
        15'h073B: data = 12'h081;
        15'h073C: data = 12'h750;
        15'h073D: data = 12'h670;
        15'h073E: data = 12'h57E;
        15'h073F: data = 12'h4AC;
        15'h0740: data = 12'h3DA;
        15'h0741: data = 12'h31F;
        15'h0742: data = 12'h50D;
        15'h0743: data = 12'h1D4;
        15'h0744: data = 12'h13F;
        15'h0745: data = 12'h0D7;
        15'h0746: data = 12'h079;
        15'h0747: data = 12'h02D;
        15'h0748: data = 12'h799;
        15'h0749: data = 12'h77F;
        15'h074A: data = 12'h764;
        15'h074B: data = 12'h786;
        15'h074C: data = 12'h7A6;
        15'h074D: data = 12'h7E0;
        15'h074E: data = 12'h75B;
        15'h074F: data = 12'h0DE;
        15'h0750: data = 12'h149;
        15'h0751: data = 12'h1CC;
        15'h0752: data = 12'h269;
        15'h0753: data = 12'h322;
        15'h0754: data = 12'h3E1;
        15'h0755: data = 12'h4B7;
        15'h0756: data = 12'h593;
        15'h0757: data = 12'h686;
        15'h0758: data = 12'h772;
        15'h0759: data = 12'h0D1;
        15'h075A: data = 12'h1A1;
        15'h075B: data = 12'h2BB;
        15'h075C: data = 12'h3CA;
        15'h075D: data = 12'h4EC;
        15'h075E: data = 12'h600;
        15'h075F: data = 12'h722;
        15'h0760: data = 12'h472;
        15'h0761: data = 12'h50D;
        15'h0762: data = 12'h2D9;
        15'h0763: data = 12'h3F5;
        15'h0764: data = 12'h507;
        15'h0765: data = 12'h607;
        15'h0766: data = 12'h6FE;
        15'h0767: data = 12'h7F0;
        15'h0768: data = 12'h116;
        15'h0769: data = 12'h1E6;
        15'h076A: data = 12'h2B4;
        15'h076B: data = 12'h378;
        15'h076C: data = 12'h425;
        15'h076D: data = 12'h4BC;
        15'h076E: data = 12'h545;
        15'h076F: data = 12'h5AC;
        15'h0770: data = 12'h5F8;
        15'h0771: data = 12'h647;
        15'h0772: data = 12'h668;
        15'h0773: data = 12'h684;
        15'h0774: data = 12'h685;
        15'h0775: data = 12'h669;
        15'h0776: data = 12'h64B;
        15'h0777: data = 12'h60F;
        15'h0778: data = 12'h5C6;
        15'h0779: data = 12'h55F;
        15'h077A: data = 12'h4E2;
        15'h077B: data = 12'h456;
        15'h077C: data = 12'h3A2;
        15'h077D: data = 12'h2E6;
        15'h077E: data = 12'h21B;
        15'h077F: data = 12'h147;
        15'h0780: data = 12'h50D;
        15'h0781: data = 12'h73A;
        15'h0782: data = 12'h642;
        15'h0783: data = 12'h542;
        15'h0784: data = 12'h42F;
        15'h0785: data = 12'h325;
        15'h0786: data = 12'h207;
        15'h0787: data = 12'h0E6;
        15'h0788: data = 12'h769;
        15'h0789: data = 12'h653;
        15'h078A: data = 12'h52F;
        15'h078B: data = 12'h415;
        15'h078C: data = 12'h2F9;
        15'h078D: data = 12'h1DB;
        15'h078E: data = 12'h0D6;
        15'h078F: data = 12'h7AC;
        15'h0790: data = 12'h6B3;
        15'h0791: data = 12'h5CA;
        15'h0792: data = 12'h4F8;
        15'h0793: data = 12'h41F;
        15'h0794: data = 12'h35D;
        15'h0795: data = 12'h2A5;
        15'h0796: data = 12'h201;
        15'h0797: data = 12'h16F;
        15'h0798: data = 12'h0F7;
        15'h0799: data = 12'h093;
        15'h079A: data = 12'h032;
        15'h079B: data = 12'h793;
        15'h079C: data = 12'h77D;
        15'h079D: data = 12'h762;
        15'h079E: data = 12'h784;
        15'h079F: data = 12'h50D;
        15'h07A0: data = 12'h7C2;
        15'h07A1: data = 12'h7FF;
        15'h07A2: data = 12'h0BB;
        15'h07A3: data = 12'h11A;
        15'h07A4: data = 12'h1A3;
        15'h07A5: data = 12'h238;
        15'h07A6: data = 12'h2E4;
        15'h07A7: data = 12'h39B;
        15'h07A8: data = 12'h46E;
        15'h07A9: data = 12'h546;
        15'h07AA: data = 12'h62F;
        15'h07AB: data = 12'h721;
        15'h07AC: data = 12'h821;
        15'h07AD: data = 12'h155;
        15'h07AE: data = 12'h25C;
        15'h07AF: data = 12'h372;
        15'h07B0: data = 12'h489;
        15'h07B1: data = 12'h59F;
        15'h07B2: data = 12'h6C9;
        15'h07B3: data = 12'h7E7;
        15'h07B4: data = 12'h159;
        15'h07B5: data = 12'h27D;
        15'h07B6: data = 12'h395;
        15'h07B7: data = 12'h4AD;
        15'h07B8: data = 12'h5B0;
        15'h07B9: data = 12'h6B7;
        15'h07BA: data = 12'h7A3;
        15'h07BB: data = 12'h0C8;
        15'h07BC: data = 12'h1A8;
        15'h07BD: data = 12'h276;
        15'h07BE: data = 12'h50D;
        15'h07BF: data = 12'h3F5;
        15'h07C0: data = 12'h494;
        15'h07C1: data = 12'h51F;
        15'h07C2: data = 12'h588;
        15'h07C3: data = 12'h5F2;
        15'h07C4: data = 12'h630;
        15'h07C5: data = 12'h66B;
        15'h07C6: data = 12'h683;
        15'h07C7: data = 12'h684;
        15'h07C8: data = 12'h685;
        15'h07C9: data = 12'h668;
        15'h07CA: data = 12'h633;
        15'h07CB: data = 12'h5E1;
        15'h07CC: data = 12'h57A;
        15'h07CD: data = 12'h50F;
        15'h07CE: data = 12'h484;
        15'h07CF: data = 12'h3E7;
        15'h07D0: data = 12'h331;
        15'h07D1: data = 12'h267;
        15'h07D2: data = 12'h18F;
        15'h07D3: data = 12'h0B1;
        15'h07D4: data = 12'h789;
        15'h07D5: data = 12'h694;
        15'h07D6: data = 12'h593;
        15'h07D7: data = 12'h496;
        15'h07D8: data = 12'h379;
        15'h07D9: data = 12'h260;
        15'h07DA: data = 12'h146;
        15'h07DB: data = 12'h023;
        15'h07DC: data = 12'h6B7;
        15'h07DD: data = 12'h50D;
        15'h07DE: data = 12'h472;
        15'h07DF: data = 12'h351;
        15'h07E0: data = 12'h23C;
        15'h07E1: data = 12'h126;
        15'h07E2: data = 12'h02D;
        15'h07E3: data = 12'h6FD;
        15'h07E4: data = 12'h614;
        15'h07E5: data = 12'h536;
        15'h07E6: data = 12'h46B;
        15'h07E7: data = 12'h39E;
        15'h07E8: data = 12'h2E3;
        15'h07E9: data = 12'h23C;
        15'h07EA: data = 12'h1A3;
        15'h07EB: data = 12'h10F;
        15'h07EC: data = 12'h0B7;
        15'h07ED: data = 12'h057;
        15'h07EE: data = 12'h7BB;
        15'h07EF: data = 12'h777;
        15'h07F0: data = 12'h776;
        15'h07F1: data = 12'h75E;
        15'h07F2: data = 12'h786;
        15'h07F3: data = 12'h7A8;
        15'h07F4: data = 12'h7E9;
        15'h07F5: data = 12'h09A;
        15'h07F6: data = 12'h0FF;
        15'h07F7: data = 12'h16D;
        15'h07F8: data = 12'h1FC;
        15'h07F9: data = 12'h29E;
        15'h07FA: data = 12'h35B;
        15'h07FB: data = 12'h428;
        15'h07FC: data = 12'h50D;
        15'h07FD: data = 12'h5E7;
        15'h07FE: data = 12'h6D7;
        15'h07FF: data = 12'h7C8;
        15'h0800: data = 12'h0FB;
        15'h0801: data = 12'h202;
        15'h0802: data = 12'h30B;
        15'h0803: data = 12'h42D;
        15'h0804: data = 12'h53D;
        15'h0805: data = 12'h663;
        15'h0806: data = 12'h78C;
        15'h0807: data = 12'h100;
        15'h0808: data = 12'h21F;
        15'h0809: data = 12'h33C;
        15'h080A: data = 12'h44E;
        15'h080B: data = 12'h55E;
        15'h080C: data = 12'h65D;
        15'h080D: data = 12'h750;
        15'h080E: data = 12'h3AE;
        15'h080F: data = 12'h160;
        15'h0810: data = 12'h235;
        15'h0811: data = 12'h2FB;
        15'h0812: data = 12'h3B6;
        15'h0813: data = 12'h45E;
        15'h0814: data = 12'h4EF;
        15'h0815: data = 12'h564;
        15'h0816: data = 12'h5D5;
        15'h0817: data = 12'h60E;
        15'h0818: data = 12'h64D;
        15'h0819: data = 12'h676;
        15'h081A: data = 12'h684;
        15'h081B: data = 12'h50D;
        15'h081C: data = 12'h668;
        15'h081D: data = 12'h63F;
        15'h081E: data = 12'h5F7;
        15'h081F: data = 12'h5A7;
        15'h0820: data = 12'h539;
        15'h0821: data = 12'h4B1;
        15'h0822: data = 12'h419;
        15'h0823: data = 12'h367;
        15'h0824: data = 12'h2AA;
        15'h0825: data = 12'h1DA;
        15'h0826: data = 12'h102;
        15'h0827: data = 12'h03E;
        15'h0828: data = 12'h6E7;
        15'h0829: data = 12'h5EC;
        15'h082A: data = 12'h4E5;
        15'h082B: data = 12'h3DA;
        15'h082C: data = 12'h2BD;
        15'h082D: data = 12'h1A3;
        15'h082E: data = 12'h082;
        15'h082F: data = 12'h70C;
        15'h0830: data = 12'h5F3;
        15'h0831: data = 12'h4D3;
        15'h0832: data = 12'h3AE;
        15'h0833: data = 12'h298;
        15'h0834: data = 12'h17F;
        15'h0835: data = 12'h086;
        15'h0836: data = 12'h74F;
        15'h0837: data = 12'h66C;
        15'h0838: data = 12'h57F;
        15'h0839: data = 12'h4A9;
        15'h083A: data = 12'h50D;
        15'h083B: data = 12'h31E;
        15'h083C: data = 12'h277;
        15'h083D: data = 12'h1D6;
        15'h083E: data = 12'h141;
        15'h083F: data = 12'h0DB;
        15'h0840: data = 12'h079;
        15'h0841: data = 12'h028;
        15'h0842: data = 12'h795;
        15'h0843: data = 12'h77A;
        15'h0844: data = 12'h75F;
        15'h0845: data = 12'h784;
        15'h0846: data = 12'h7AA;
        15'h0847: data = 12'h7E3;
        15'h0848: data = 12'h703;
        15'h0849: data = 12'h0DC;
        15'h084A: data = 12'h144;
        15'h084B: data = 12'h1C8;
        15'h084C: data = 12'h267;
        15'h084D: data = 12'h31F;
        15'h084E: data = 12'h3E3;
        15'h084F: data = 12'h4B5;
        15'h0850: data = 12'h595;
        15'h0851: data = 12'h685;
        15'h0852: data = 12'h777;
        15'h0853: data = 12'h0CF;
        15'h0854: data = 12'h1A5;
        15'h0855: data = 12'h2BB;
        15'h0856: data = 12'h3CC;
        15'h0857: data = 12'h4F4;
        15'h0858: data = 12'h608;
        15'h0859: data = 12'h50D;
        15'h085A: data = 12'h3AC;
        15'h085B: data = 12'h1BA;
        15'h085C: data = 12'h2D9;
        15'h085D: data = 12'h3FA;
        15'h085E: data = 12'h509;
        15'h085F: data = 12'h60F;
        15'h0860: data = 12'h707;
        15'h0861: data = 12'h7F9;
        15'h0862: data = 12'h118;
        15'h0863: data = 12'h1EB;
        15'h0864: data = 12'h2B8;
        15'h0865: data = 12'h378;
        15'h0866: data = 12'h421;
        15'h0867: data = 12'h4C0;
        15'h0868: data = 12'h548;
        15'h0869: data = 12'h5B6;
        15'h086A: data = 12'h5FF;
        15'h086B: data = 12'h64C;
        15'h086C: data = 12'h66D;
        15'h086D: data = 12'h687;
        15'h086E: data = 12'h683;
        15'h086F: data = 12'h66A;
        15'h0870: data = 12'h649;
        15'h0871: data = 12'h60D;
        15'h0872: data = 12'h5C4;
        15'h0873: data = 12'h55F;
        15'h0874: data = 12'h4D9;
        15'h0875: data = 12'h451;
        15'h0876: data = 12'h3A7;
        15'h0877: data = 12'h2EE;
        15'h0878: data = 12'h50D;
        15'h0879: data = 12'h14A;
        15'h087A: data = 12'h069;
        15'h087B: data = 12'h739;
        15'h087C: data = 12'h63C;
        15'h087D: data = 12'h53B;
        15'h087E: data = 12'h42B;
        15'h087F: data = 12'h322;
        15'h0880: data = 12'h204;
        15'h0881: data = 12'h0EF;
        15'h0882: data = 12'h76D;
        15'h0883: data = 12'h659;
        15'h0884: data = 12'h530;
        15'h0885: data = 12'h418;
        15'h0886: data = 12'h2F0;
        15'h0887: data = 12'h1DA;
        15'h0888: data = 12'h0D5;
        15'h0889: data = 12'h7AB;
        15'h088A: data = 12'h6B0;
        15'h088B: data = 12'h5CB;
        15'h088C: data = 12'h4F9;
        15'h088D: data = 12'h41E;
        15'h088E: data = 12'h35A;
        15'h088F: data = 12'h2A7;
        15'h0890: data = 12'h203;
        15'h0891: data = 12'h176;
        15'h0892: data = 12'h102;
        15'h0893: data = 12'h097;
        15'h0894: data = 12'h03A;
        15'h0895: data = 12'h793;
        15'h0896: data = 12'h776;
        15'h0897: data = 12'h50D;
        15'h0898: data = 12'h77F;
        15'h0899: data = 12'h781;
        15'h089A: data = 12'h7C4;
        15'h089B: data = 12'h804;
        15'h089C: data = 12'h0C3;
        15'h089D: data = 12'h122;
        15'h089E: data = 12'h1A8;
        15'h089F: data = 12'h237;
        15'h08A0: data = 12'h2E1;
        15'h08A1: data = 12'h39A;
        15'h08A2: data = 12'h46D;
        15'h08A3: data = 12'h544;
        15'h08A4: data = 12'h632;
        15'h08A5: data = 12'h723;
        15'h08A6: data = 12'h81E;
        15'h08A7: data = 12'h155;
        15'h08A8: data = 12'h261;
        15'h08A9: data = 12'h37A;
        15'h08AA: data = 12'h48A;
        15'h08AB: data = 12'h5A1;
        15'h08AC: data = 12'h6CA;
        15'h08AD: data = 12'h7E7;
        15'h08AE: data = 12'h153;
        15'h08AF: data = 12'h27D;
        15'h08B0: data = 12'h396;
        15'h08B1: data = 12'h4AC;
        15'h08B2: data = 12'h5B5;
        15'h08B3: data = 12'h6C0;
        15'h08B4: data = 12'h7A9;
        15'h08B5: data = 12'h0D2;
        15'h08B6: data = 12'h50D;
        15'h08B7: data = 12'h279;
        15'h08B8: data = 12'h333;
        15'h08B9: data = 12'h3EE;
        15'h08BA: data = 12'h495;
        15'h08BB: data = 12'h518;
        15'h08BC: data = 12'h58C;
        15'h08BD: data = 12'h5F6;
        15'h08BE: data = 12'h637;
        15'h08BF: data = 12'h674;
        15'h08C0: data = 12'h68F;
        15'h08C1: data = 12'h68B;
        15'h08C2: data = 12'h688;
        15'h08C3: data = 12'h664;
        15'h08C4: data = 12'h628;
        15'h08C5: data = 12'h5DC;
        15'h08C6: data = 12'h573;
        15'h08C7: data = 12'h511;
        15'h08C8: data = 12'h483;
        15'h08C9: data = 12'h3E5;
        15'h08CA: data = 12'h336;
        15'h08CB: data = 12'h272;
        15'h08CC: data = 12'h197;
        15'h08CD: data = 12'h0BA;
        15'h08CE: data = 12'h78E;
        15'h08CF: data = 12'h692;
        15'h08D0: data = 12'h58E;
        15'h08D1: data = 12'h486;
        15'h08D2: data = 12'h36E;
        15'h08D3: data = 12'h261;
        15'h08D4: data = 12'h149;
        15'h08D5: data = 12'h50D;
        15'h08D6: data = 12'h6BB;
        15'h08D7: data = 12'h593;
        15'h08D8: data = 12'h47D;
        15'h08D9: data = 12'h357;
        15'h08DA: data = 12'h23A;
        15'h08DB: data = 12'h124;
        15'h08DC: data = 12'h027;
        15'h08DD: data = 12'h6F8;
        15'h08DE: data = 12'h60D;
        15'h08DF: data = 12'h52D;
        15'h08E0: data = 12'h465;
        15'h08E1: data = 12'h39B;
        15'h08E2: data = 12'h2E4;
        15'h08E3: data = 12'h23F;
        15'h08E4: data = 12'h1A9;
        15'h08E5: data = 12'h11E;
        15'h08E6: data = 12'h0BF;
        15'h08E7: data = 12'h05A;
        15'h08E8: data = 12'h79D;
        15'h08E9: data = 12'h773;
        15'h08EA: data = 12'h76C;
        15'h08EB: data = 12'h756;
        15'h08EC: data = 12'h779;
        15'h08ED: data = 12'h7A2;
        15'h08EE: data = 12'h7E8;
        15'h08EF: data = 12'h0A1;
        15'h08F0: data = 12'h109;
        15'h08F1: data = 12'h179;
        15'h08F2: data = 12'h20D;
        15'h08F3: data = 12'h2AB;
        15'h08F4: data = 12'h50D;
        15'h08F5: data = 12'h422;
        15'h08F6: data = 12'h4F5;
        15'h08F7: data = 12'h5DA;
        15'h08F8: data = 12'h6D0;
        15'h08F9: data = 12'h7CB;
        15'h08FA: data = 12'h104;
        15'h08FB: data = 12'h20A;
        15'h08FC: data = 12'h31A;
        15'h08FD: data = 12'h437;
        15'h08FE: data = 12'h543;
        15'h08FF: data = 12'h65F;
        15'h0900: data = 12'h785;
        15'h0901: data = 12'h0EB;
        15'h0902: data = 12'h20D;
        15'h0903: data = 12'h336;
        15'h0904: data = 12'h44A;
        15'h0905: data = 12'h560;
        15'h0906: data = 12'h662;
        15'h0907: data = 12'h75C;
        15'h0908: data = 12'h55E;
        15'h0909: data = 12'h162;
        15'h090A: data = 12'h232;
        15'h090B: data = 12'h2F6;
        15'h090C: data = 12'h3AB;
        15'h090D: data = 12'h450;
        15'h090E: data = 12'h4E6;
        15'h090F: data = 12'h55D;
        15'h0910: data = 12'h5D3;
        15'h0911: data = 12'h61C;
        15'h0912: data = 12'h658;
        15'h0913: data = 12'h50D;
        15'h0914: data = 12'h68F;
        15'h0915: data = 12'h689;
        15'h0916: data = 12'h667;
        15'h0917: data = 12'h635;
        15'h0918: data = 12'h5E4;
        15'h0919: data = 12'h596;
        15'h091A: data = 12'h537;
        15'h091B: data = 12'h4B1;
        15'h091C: data = 12'h419;
        15'h091D: data = 12'h372;
        15'h091E: data = 12'h2B6;
        15'h091F: data = 12'h1E5;
        15'h0920: data = 12'h10F;
        15'h0921: data = 12'h01C;
        15'h0922: data = 12'h6E4;
        15'h0923: data = 12'h5E8;
        15'h0924: data = 12'h4DC;
        15'h0925: data = 12'h3D0;
        15'h0926: data = 12'h2B4;
        15'h0927: data = 12'h1A0;
        15'h0928: data = 12'h087;
        15'h0929: data = 12'h70F;
        15'h092A: data = 12'h5F7;
        15'h092B: data = 12'h4E2;
        15'h092C: data = 12'h3BC;
        15'h092D: data = 12'h2AA;
        15'h092E: data = 12'h18D;
        15'h092F: data = 12'h086;
        15'h0930: data = 12'h746;
        15'h0931: data = 12'h65D;
        15'h0932: data = 12'h50D;
        15'h0933: data = 12'h49E;
        15'h0934: data = 12'h3D3;
        15'h0935: data = 12'h31A;
        15'h0936: data = 12'h276;
        15'h0937: data = 12'h1DD;
        15'h0938: data = 12'h14B;
        15'h0939: data = 12'h0E6;
        15'h093A: data = 12'h080;
        15'h093B: data = 12'h02E;
        15'h093C: data = 12'h795;
        15'h093D: data = 12'h770;
        15'h093E: data = 12'h755;
        15'h093F: data = 12'h774;
        15'h0940: data = 12'h799;
        15'h0941: data = 12'h7DB;
        15'h0942: data = 12'h81F;
        15'h0943: data = 12'h0E3;
        15'h0944: data = 12'h153;
        15'h0945: data = 12'h1E1;
        15'h0946: data = 12'h277;
        15'h0947: data = 12'h328;
        15'h0948: data = 12'h3E0;
        15'h0949: data = 12'h4AC;
        15'h094A: data = 12'h586;
        15'h094B: data = 12'h675;
        15'h094C: data = 12'h76B;
        15'h094D: data = 12'h0E0;
        15'h094E: data = 12'h1A7;
        15'h094F: data = 12'h2C9;
        15'h0950: data = 12'h3DC;
        15'h0951: data = 12'h50D;
        15'h0952: data = 12'h60D;
        15'h0953: data = 12'h71D;
        15'h0954: data = 12'h40C;
        15'h0955: data = 12'h1AD;
        15'h0956: data = 12'h2CD;
        15'h0957: data = 12'h3EC;
        15'h0958: data = 12'h506;
        15'h0959: data = 12'h614;
        15'h095A: data = 12'h70F;
        15'h095B: data = 12'h800;
        15'h095C: data = 12'h121;
        15'h095D: data = 12'h1F1;
        15'h095E: data = 12'h2B5;
        15'h095F: data = 12'h370;
        15'h0960: data = 12'h411;
        15'h0961: data = 12'h4AF;
        15'h0962: data = 12'h539;
        15'h0963: data = 12'h5AB;
        15'h0964: data = 12'h5F5;
        15'h0965: data = 12'h64F;
        15'h0966: data = 12'h675;
        15'h0967: data = 12'h696;
        15'h0968: data = 12'h693;
        15'h0969: data = 12'h66E;
        15'h096A: data = 12'h64C;
        15'h096B: data = 12'h604;
        15'h096C: data = 12'h5B9;
        15'h096D: data = 12'h54B;
        15'h096E: data = 12'h4D5;
        15'h096F: data = 12'h452;
        15'h0970: data = 12'h50D;
        15'h0971: data = 12'h2F8;
        15'h0972: data = 12'h22B;
        15'h0973: data = 12'h155;
        15'h0974: data = 12'h077;
        15'h0975: data = 12'h744;
        15'h0976: data = 12'h643;
        15'h0977: data = 12'h539;
        15'h0978: data = 12'h422;
        15'h0979: data = 12'h312;
        15'h097A: data = 12'h1F2;
        15'h097B: data = 12'h0DC;
        15'h097C: data = 12'h77A;
        15'h097D: data = 12'h659;
        15'h097E: data = 12'h537;
        15'h097F: data = 12'h422;
        15'h0980: data = 12'h302;
        15'h0981: data = 12'h1EC;
        15'h0982: data = 12'h0DE;
        15'h0983: data = 12'h794;
        15'h0984: data = 12'h6AC;
        15'h0985: data = 12'h5BF;
        15'h0986: data = 12'h4E3;
        15'h0987: data = 12'h410;
        15'h0988: data = 12'h34C;
        15'h0989: data = 12'h29C;
        15'h098A: data = 12'h1FF;
        15'h098B: data = 12'h17A;
        15'h098C: data = 12'h10D;
        15'h098D: data = 12'h0A9;
        15'h098E: data = 12'h04B;
        15'h098F: data = 12'h50D;
        15'h0990: data = 12'h77A;
        15'h0991: data = 12'h754;
        15'h0992: data = 12'h774;
        15'h0993: data = 12'h771;
        15'h0994: data = 12'h7B6;
        15'h0995: data = 12'h7F6;
        15'h0996: data = 12'h0BF;
        15'h0997: data = 12'h125;
        15'h0998: data = 12'h1BB;
        15'h0999: data = 12'h24A;
        15'h099A: data = 12'h2F6;
        15'h099B: data = 12'h3AB;
        15'h099C: data = 12'h474;
        15'h099D: data = 12'h53D;
        15'h099E: data = 12'h628;
        15'h099F: data = 12'h710;
        15'h09A0: data = 12'h815;
        15'h09A1: data = 12'h14C;
        15'h09A2: data = 12'h25F;
        15'h09A3: data = 12'h382;
        15'h09A4: data = 12'h498;
        15'h09A5: data = 12'h5AE;
        15'h09A6: data = 12'h6D8;
        15'h09A7: data = 12'h7E9;
        15'h09A8: data = 12'h153;
        15'h09A9: data = 12'h272;
        15'h09AA: data = 12'h385;
        15'h09AB: data = 12'h4A1;
        15'h09AC: data = 12'h5AC;
        15'h09AD: data = 12'h6BD;
        15'h09AE: data = 12'h50D;
        15'h09AF: data = 12'h0DD;
        15'h09B0: data = 12'h1BB;
        15'h09B1: data = 12'h28A;
        15'h09B2: data = 12'h33C;
        15'h09B3: data = 12'h3EB;
        15'h09B4: data = 12'h488;
        15'h09B5: data = 12'h50F;
        15'h09B6: data = 12'h578;
        15'h09B7: data = 12'h5E8;
        15'h09B8: data = 12'h635;
        15'h09B9: data = 12'h677;
        15'h09BA: data = 12'h695;
        15'h09BB: data = 12'h698;
        15'h09BC: data = 12'h693;
        15'h09BD: data = 12'h66A;
        15'h09BE: data = 12'h627;
        15'h09BF: data = 12'h5CF;
        15'h09C0: data = 12'h564;
        15'h09C1: data = 12'h4FB;
        15'h09C2: data = 12'h472;
        15'h09C3: data = 12'h3DE;
        15'h09C4: data = 12'h32F;
        15'h09C5: data = 12'h272;
        15'h09C6: data = 12'h19C;
        15'h09C7: data = 12'h0C3;
        15'h09C8: data = 12'h78A;
        15'h09C9: data = 12'h6A0;
        15'h09CA: data = 12'h599;
        15'h09CB: data = 12'h48C;
        15'h09CC: data = 12'h36C;
        15'h09CD: data = 12'h50D;
        15'h09CE: data = 12'h135;
        15'h09CF: data = 12'h055;
        15'h09D0: data = 12'h6AB;
        15'h09D1: data = 12'h589;
        15'h09D2: data = 12'h47D;
        15'h09D3: data = 12'h361;
        15'h09D4: data = 12'h24B;
        15'h09D5: data = 12'h136;
        15'h09D6: data = 12'h036;
        15'h09D7: data = 12'h706;
        15'h09D8: data = 12'h610;
        15'h09D9: data = 12'h529;
        15'h09DA: data = 12'h45C;
        15'h09DB: data = 12'h38B;
        15'h09DC: data = 12'h2D4;
        15'h09DD: data = 12'h22D;
        15'h09DE: data = 12'h19E;
        15'h09DF: data = 12'h11C;
        15'h09E0: data = 12'h0C8;
        15'h09E1: data = 12'h067;
        15'h09E2: data = 12'h75A;
        15'h09E3: data = 12'h782;
        15'h09E4: data = 12'h779;
        15'h09E5: data = 12'h75E;
        15'h09E6: data = 12'h779;
        15'h09E7: data = 12'h797;
        15'h09E8: data = 12'h7DB;
        15'h09E9: data = 12'h091;
        15'h09EA: data = 12'h0FC;
        15'h09EB: data = 12'h178;
        15'h09EC: data = 12'h50D;
        15'h09ED: data = 12'h2BB;
        15'h09EE: data = 12'h36E;
        15'h09EF: data = 12'h433;
        15'h09F0: data = 12'h502;
        15'h09F1: data = 12'h5E4;
        15'h09F2: data = 12'h6C9;
        15'h09F3: data = 12'h7BD;
        15'h09F4: data = 12'h0F1;
        15'h09F5: data = 12'h1FF;
        15'h09F6: data = 12'h313;
        15'h09F7: data = 12'h43C;
        15'h09F8: data = 12'h553;
        15'h09F9: data = 12'h673;
        15'h09FA: data = 12'h797;
        15'h09FB: data = 12'h0FB;
        15'h09FC: data = 12'h215;
        15'h09FD: data = 12'h333;
        15'h09FE: data = 12'h449;
        15'h09FF: data = 12'h558;
        15'h0A00: data = 12'h65A;
        15'h0A01: data = 12'h759;
        15'h0A02: data = 12'h1EC;
        15'h0A03: data = 12'h173;
        15'h0A04: data = 12'h243;
        15'h0A05: data = 12'h304;
        15'h0A06: data = 12'h3BD;
        15'h0A07: data = 12'h457;
        15'h0A08: data = 12'h4E5;
        15'h0A09: data = 12'h551;
        15'h0A0A: data = 12'h5C6;
        15'h0A0B: data = 12'h50D;
        15'h0A0C: data = 12'h64C;
        15'h0A0D: data = 12'h688;
        15'h0A0E: data = 12'h698;
        15'h0A0F: data = 12'h69E;
        15'h0A10: data = 12'h67A;
        15'h0A11: data = 12'h641;
        15'h0A12: data = 12'h5F1;
        15'h0A13: data = 12'h597;
        15'h0A14: data = 12'h52D;
        15'h0A15: data = 12'h49F;
        15'h0A16: data = 12'h411;
        15'h0A17: data = 12'h362;
        15'h0A18: data = 12'h2A9;
        15'h0A19: data = 12'h1DF;
        15'h0A1A: data = 12'h10A;
        15'h0A1B: data = 12'h0C8;
        15'h0A1C: data = 12'h6F6;
        15'h0A1D: data = 12'h5FB;
        15'h0A1E: data = 12'h4F0;
        15'h0A1F: data = 12'h3DA;
        15'h0A20: data = 12'h2B6;
        15'h0A21: data = 12'h196;
        15'h0A22: data = 12'h076;
        15'h0A23: data = 12'h6F8;
        15'h0A24: data = 12'h5E5;
        15'h0A25: data = 12'h4D2;
        15'h0A26: data = 12'h3B0;
        15'h0A27: data = 12'h2A3;
        15'h0A28: data = 12'h194;
        15'h0A29: data = 12'h093;
        15'h0A2A: data = 12'h50D;
        15'h0A2B: data = 12'h670;
        15'h0A2C: data = 12'h57C;
        15'h0A2D: data = 12'h4A3;
        15'h0A2E: data = 12'h3CE;
        15'h0A2F: data = 12'h310;
        15'h0A30: data = 12'h262;
        15'h0A31: data = 12'h1CA;
        15'h0A32: data = 12'h13C;
        15'h0A33: data = 12'h0DC;
        15'h0A34: data = 12'h085;
        15'h0A35: data = 12'h03A;
        15'h0A36: data = 12'h7A9;
        15'h0A37: data = 12'h787;
        15'h0A38: data = 12'h765;
        15'h0A39: data = 12'h784;
        15'h0A3A: data = 12'h79A;
        15'h0A3B: data = 12'h7CE;
        15'h0A3C: data = 12'h53E;
        15'h0A3D: data = 12'h0D1;
        15'h0A3E: data = 12'h144;
        15'h0A3F: data = 12'h1CF;
        15'h0A40: data = 12'h277;
        15'h0A41: data = 12'h333;
        15'h0A42: data = 12'h3F0;
        15'h0A43: data = 12'h4BA;
        15'h0A44: data = 12'h597;
        15'h0A45: data = 12'h680;
        15'h0A46: data = 12'h76F;
        15'h0A47: data = 12'h1AA;
        15'h0A48: data = 12'h198;
        15'h0A49: data = 12'h50D;
        15'h0A4A: data = 12'h3CB;
        15'h0A4B: data = 12'h4F0;
        15'h0A4C: data = 12'h613;
        15'h0A4D: data = 12'h729;
        15'h0A4E: data = 12'h724;
        15'h0A4F: data = 12'h1BC;
        15'h0A50: data = 12'h2D7;
        15'h0A51: data = 12'h3F0;
        15'h0A52: data = 12'h4FE;
        15'h0A53: data = 12'h603;
        15'h0A54: data = 12'h6FD;
        15'h0A55: data = 12'h7F4;
        15'h0A56: data = 12'h11F;
        15'h0A57: data = 12'h1F2;
        15'h0A58: data = 12'h2C0;
        15'h0A59: data = 12'h37D;
        15'h0A5A: data = 12'h427;
        15'h0A5B: data = 12'h4B9;
        15'h0A5C: data = 12'h53F;
        15'h0A5D: data = 12'h5A4;
        15'h0A5E: data = 12'h5EB;
        15'h0A5F: data = 12'h644;
        15'h0A60: data = 12'h665;
        15'h0A61: data = 12'h686;
        15'h0A62: data = 12'h68A;
        15'h0A63: data = 12'h676;
        15'h0A64: data = 12'h655;
        15'h0A65: data = 12'h616;
        15'h0A66: data = 12'h5C7;
        15'h0A67: data = 12'h559;
        15'h0A68: data = 12'h50D;
        15'h0A69: data = 12'h447;
        15'h0A6A: data = 12'h39A;
        15'h0A6B: data = 12'h2E8;
        15'h0A6C: data = 12'h21B;
        15'h0A6D: data = 12'h147;
        15'h0A6E: data = 12'h068;
        15'h0A6F: data = 12'h73C;
        15'h0A70: data = 12'h645;
        15'h0A71: data = 12'h545;
        15'h0A72: data = 12'h432;
        15'h0A73: data = 12'h321;
        15'h0A74: data = 12'h203;
        15'h0A75: data = 12'h0E9;
        15'h0A76: data = 12'h76F;
        15'h0A77: data = 12'h64C;
        15'h0A78: data = 12'h525;
        15'h0A79: data = 12'h40E;
        15'h0A7A: data = 12'h2F6;
        15'h0A7B: data = 12'h1DD;
        15'h0A7C: data = 12'h0DC;
        15'h0A7D: data = 12'h7B5;
        15'h0A7E: data = 12'h6BA;
        15'h0A7F: data = 12'h5CF;
        15'h0A80: data = 12'h4F6;
        15'h0A81: data = 12'h41F;
        15'h0A82: data = 12'h358;
        15'h0A83: data = 12'h2A1;
        15'h0A84: data = 12'h1F7;
        15'h0A85: data = 12'h16C;
        15'h0A86: data = 12'h0F4;
        15'h0A87: data = 12'h50D;
        15'h0A88: data = 12'h036;
        15'h0A89: data = 12'h798;
        15'h0A8A: data = 12'h780;
        15'h0A8B: data = 12'h763;
        15'h0A8C: data = 12'h781;
        15'h0A8D: data = 12'h785;
        15'h0A8E: data = 12'h7BC;
        15'h0A8F: data = 12'h802;
        15'h0A90: data = 12'h0BA;
        15'h0A91: data = 12'h11B;
        15'h0A92: data = 12'h1A4;
        15'h0A93: data = 12'h23B;
        15'h0A94: data = 12'h2E1;
        15'h0A95: data = 12'h3A0;
        15'h0A96: data = 12'h473;
        15'h0A97: data = 12'h54A;
        15'h0A98: data = 12'h634;
        15'h0A99: data = 12'h725;
        15'h0A9A: data = 12'h823;
        15'h0A9B: data = 12'h152;
        15'h0A9C: data = 12'h259;
        15'h0A9D: data = 12'h36D;
        15'h0A9E: data = 12'h486;
        15'h0A9F: data = 12'h59E;
        15'h0AA0: data = 12'h6CB;
        15'h0AA1: data = 12'h7EC;
        15'h0AA2: data = 12'h15B;
        15'h0AA3: data = 12'h283;
        15'h0AA4: data = 12'h399;
        15'h0AA5: data = 12'h4B0;
        15'h0AA6: data = 12'h50D;
        15'h0AA7: data = 12'h6B4;
        15'h0AA8: data = 12'h79F;
        15'h0AA9: data = 12'h0D2;
        15'h0AAA: data = 12'h1AA;
        15'h0AAB: data = 12'h27C;
        15'h0AAC: data = 12'h33B;
        15'h0AAD: data = 12'h3F4;
        15'h0AAE: data = 12'h498;
        15'h0AAF: data = 12'h51E;
        15'h0AB0: data = 12'h58A;
        15'h0AB1: data = 12'h5F1;
        15'h0AB2: data = 12'h62F;
        15'h0AB3: data = 12'h668;
        15'h0AB4: data = 12'h685;
        15'h0AB5: data = 12'h686;
        15'h0AB6: data = 12'h689;
        15'h0AB7: data = 12'h665;
        15'h0AB8: data = 12'h631;
        15'h0AB9: data = 12'h5DF;
        15'h0ABA: data = 12'h576;
        15'h0ABB: data = 12'h50D;
        15'h0ABC: data = 12'h483;
        15'h0ABD: data = 12'h3E3;
        15'h0ABE: data = 12'h330;
        15'h0ABF: data = 12'h267;
        15'h0AC0: data = 12'h18E;
        15'h0AC1: data = 12'h0AE;
        15'h0AC2: data = 12'h78B;
        15'h0AC3: data = 12'h694;
        15'h0AC4: data = 12'h592;
        15'h0AC5: data = 12'h50D;
        15'h0AC6: data = 12'h37B;
        15'h0AC7: data = 12'h260;
        15'h0AC8: data = 12'h147;
        15'h0AC9: data = 12'h023;
        15'h0ACA: data = 12'h6B6;
        15'h0ACB: data = 12'h58B;
        15'h0ACC: data = 12'h472;
        15'h0ACD: data = 12'h352;
        15'h0ACE: data = 12'h23C;
        15'h0ACF: data = 12'h12A;
        15'h0AD0: data = 12'h02D;
        15'h0AD1: data = 12'h6FC;
        15'h0AD2: data = 12'h611;
        15'h0AD3: data = 12'h530;
        15'h0AD4: data = 12'h467;
        15'h0AD5: data = 12'h39A;
        15'h0AD6: data = 12'h2E1;
        15'h0AD7: data = 12'h237;
        15'h0AD8: data = 12'h19A;
        15'h0AD9: data = 12'h10F;
        15'h0ADA: data = 12'h0B6;
        15'h0ADB: data = 12'h054;
        15'h0ADC: data = 12'h7B0;
        15'h0ADD: data = 12'h774;
        15'h0ADE: data = 12'h770;
        15'h0ADF: data = 12'h763;
        15'h0AE0: data = 12'h786;
        15'h0AE1: data = 12'h7A6;
        15'h0AE2: data = 12'h7ED;
        15'h0AE3: data = 12'h09A;
        15'h0AE4: data = 12'h50D;
        15'h0AE5: data = 12'h173;
        15'h0AE6: data = 12'h202;
        15'h0AE7: data = 12'h2A2;
        15'h0AE8: data = 12'h35C;
        15'h0AE9: data = 12'h428;
        15'h0AEA: data = 12'h502;
        15'h0AEB: data = 12'h5EA;
        15'h0AEC: data = 12'h6DA;
        15'h0AED: data = 12'h7CE;
        15'h0AEE: data = 12'h103;
        15'h0AEF: data = 12'h207;
        15'h0AF0: data = 12'h30E;
        15'h0AF1: data = 12'h42C;
        15'h0AF2: data = 12'h53D;
        15'h0AF3: data = 12'h661;
        15'h0AF4: data = 12'h788;
        15'h0AF5: data = 12'h0FB;
        15'h0AF6: data = 12'h21D;
        15'h0AF7: data = 12'h337;
        15'h0AF8: data = 12'h455;
        15'h0AF9: data = 12'h55D;
        15'h0AFA: data = 12'h65F;
        15'h0AFB: data = 12'h756;
        15'h0AFC: data = 12'h3FF;
        15'h0AFD: data = 12'h166;
        15'h0AFE: data = 12'h234;
        15'h0AFF: data = 12'h2F9;
        15'h0B00: data = 12'h3B1;
        15'h0B01: data = 12'h45C;
        15'h0B02: data = 12'h4F3;
        15'h0B03: data = 12'h50D;
        15'h0B04: data = 12'h5D2;
        15'h0B05: data = 12'h615;
        15'h0B06: data = 12'h657;
        15'h0B07: data = 12'h67B;
        15'h0B08: data = 12'h684;
        15'h0B09: data = 12'h687;
        15'h0B0A: data = 12'h663;
        15'h0B0B: data = 12'h636;
        15'h0B0C: data = 12'h5EB;
        15'h0B0D: data = 12'h5A0;
        15'h0B0E: data = 12'h53C;
        15'h0B0F: data = 12'h4B0;
        15'h0B10: data = 12'h419;
        15'h0B11: data = 12'h36A;
        15'h0B12: data = 12'h2AD;
        15'h0B13: data = 12'h1D9;
        15'h0B14: data = 12'h0FE;
        15'h0B15: data = 12'h022;
        15'h0B16: data = 12'h6E4;
        15'h0B17: data = 12'h5EB;
        15'h0B18: data = 12'h4E2;
        15'h0B19: data = 12'h3D9;
        15'h0B1A: data = 12'h2BF;
        15'h0B1B: data = 12'h1A6;
        15'h0B1C: data = 12'h087;
        15'h0B1D: data = 12'h70A;
        15'h0B1E: data = 12'h5F4;
        15'h0B1F: data = 12'h4D9;
        15'h0B20: data = 12'h3AF;
        15'h0B21: data = 12'h29B;
        15'h0B22: data = 12'h50D;
        15'h0B23: data = 12'h07F;
        15'h0B24: data = 12'h745;
        15'h0B25: data = 12'h664;
        15'h0B26: data = 12'h573;
        15'h0B27: data = 12'h4A7;
        15'h0B28: data = 12'h3DB;
        15'h0B29: data = 12'h323;
        15'h0B2A: data = 12'h278;
        15'h0B2B: data = 12'h1DB;
        15'h0B2C: data = 12'h145;
        15'h0B2D: data = 12'h0DA;
        15'h0B2E: data = 12'h077;
        15'h0B2F: data = 12'h7A6;
        15'h0B30: data = 12'h791;
        15'h0B31: data = 12'h777;
        15'h0B32: data = 12'h75D;
        15'h0B33: data = 12'h780;
        15'h0B34: data = 12'h7A4;
        15'h0B35: data = 12'h7DC;
        15'h0B36: data = 12'h803;
        15'h0B37: data = 12'h0E0;
        15'h0B38: data = 12'h14D;
        15'h0B39: data = 12'h1D1;
        15'h0B3A: data = 12'h26D;
        15'h0B3B: data = 12'h322;
        15'h0B3C: data = 12'h3E1;
        15'h0B3D: data = 12'h4B0;
        15'h0B3E: data = 12'h58F;
        15'h0B3F: data = 12'h687;
        15'h0B40: data = 12'h774;
        15'h0B41: data = 12'h50D;
        15'h0B42: data = 12'h1A9;
        15'h0B43: data = 12'h2C2;
        15'h0B44: data = 12'h3D2;
        15'h0B45: data = 12'h4F4;
        15'h0B46: data = 12'h602;
        15'h0B47: data = 12'h720;
        15'h0B48: data = 12'h34B;
        15'h0B49: data = 12'h1B6;
        15'h0B4A: data = 12'h2DA;
        15'h0B4B: data = 12'h3FB;
        15'h0B4C: data = 12'h50B;
        15'h0B4D: data = 12'h611;
        15'h0B4E: data = 12'h70E;
        15'h0B4F: data = 12'h7F8;
        15'h0B50: data = 12'h119;
        15'h0B51: data = 12'h1EB;
        15'h0B52: data = 12'h2B7;
        15'h0B53: data = 12'h371;
        15'h0B54: data = 12'h41E;
        15'h0B55: data = 12'h4BC;
        15'h0B56: data = 12'h544;
        15'h0B57: data = 12'h5AE;
        15'h0B58: data = 12'h5FC;
        15'h0B59: data = 12'h64D;
        15'h0B5A: data = 12'h66A;
        15'h0B5B: data = 12'h687;
        15'h0B5C: data = 12'h683;
        15'h0B5D: data = 12'h667;
        15'h0B5E: data = 12'h647;
        15'h0B5F: data = 12'h609;
        15'h0B60: data = 12'h50D;
        15'h0B61: data = 12'h557;
        15'h0B62: data = 12'h4DD;
        15'h0B63: data = 12'h455;
        15'h0B64: data = 12'h3A5;
        15'h0B65: data = 12'h2F5;
        15'h0B66: data = 12'h224;
        15'h0B67: data = 12'h149;
        15'h0B68: data = 12'h063;
        15'h0B69: data = 12'h731;
        15'h0B6A: data = 12'h63A;
        15'h0B6B: data = 12'h535;
        15'h0B6C: data = 12'h427;
        15'h0B6D: data = 12'h31D;
        15'h0B6E: data = 12'h204;
        15'h0B6F: data = 12'h0E9;
        15'h0B70: data = 12'h763;
        15'h0B71: data = 12'h652;
        15'h0B72: data = 12'h532;
        15'h0B73: data = 12'h41A;
        15'h0B74: data = 12'h2F7;
        15'h0B75: data = 12'h1D9;
        15'h0B76: data = 12'h0D1;
        15'h0B77: data = 12'h7A8;
        15'h0B78: data = 12'h6AB;
        15'h0B79: data = 12'h5C7;
        15'h0B7A: data = 12'h4F3;
        15'h0B7B: data = 12'h41D;
        15'h0B7C: data = 12'h357;
        15'h0B7D: data = 12'h2A8;
        15'h0B7E: data = 12'h207;
        15'h0B7F: data = 12'h50D;
        15'h0B80: data = 12'h0FF;
        15'h0B81: data = 12'h09C;
        15'h0B82: data = 12'h03C;
        15'h0B83: data = 12'h793;
        15'h0B84: data = 12'h772;
        15'h0B85: data = 12'h754;
        15'h0B86: data = 12'h77B;
        15'h0B87: data = 12'h77D;
        15'h0B88: data = 12'h7C1;
        15'h0B89: data = 12'h801;
        15'h0B8A: data = 12'h0C6;
        15'h0B8B: data = 12'h125;
        15'h0B8C: data = 12'h1AE;
        15'h0B8D: data = 12'h23D;
        15'h0B8E: data = 12'h2E3;
        15'h0B8F: data = 12'h39C;
        15'h0B90: data = 12'h467;
        15'h0B91: data = 12'h543;
        15'h0B92: data = 12'h62E;
        15'h0B93: data = 12'h721;
        15'h0B94: data = 12'h825;
        15'h0B95: data = 12'h15C;
        15'h0B96: data = 12'h260;
        15'h0B97: data = 12'h378;
        15'h0B98: data = 12'h48D;
        15'h0B99: data = 12'h5A3;
        15'h0B9A: data = 12'h6CE;
        15'h0B9B: data = 12'h7E0;
        15'h0B9C: data = 12'h154;
        15'h0B9D: data = 12'h27D;
        15'h0B9E: data = 12'h50D;
        15'h0B9F: data = 12'h4B3;
        15'h0BA0: data = 12'h5B5;
        15'h0BA1: data = 12'h6BD;
        15'h0BA2: data = 12'h7AA;
        15'h0BA3: data = 12'h0D5;
        15'h0BA4: data = 12'h1AD;
        15'h0BA5: data = 12'h279;
        15'h0BA6: data = 12'h334;
        15'h0BA7: data = 12'h3EE;
        15'h0BA8: data = 12'h492;
        15'h0BA9: data = 12'h520;
        15'h0BAA: data = 12'h58E;
        15'h0BAB: data = 12'h5F8;
        15'h0BAC: data = 12'h636;
        15'h0BAD: data = 12'h671;
        15'h0BAE: data = 12'h689;
        15'h0BAF: data = 12'h685;
        15'h0BB0: data = 12'h683;
        15'h0BB1: data = 12'h661;
        15'h0BB2: data = 12'h628;
        15'h0BB3: data = 12'h5D9;
        15'h0BB4: data = 12'h572;
        15'h0BB5: data = 12'h50B;
        15'h0BB6: data = 12'h480;
        15'h0BB7: data = 12'h3E5;
        15'h0BB8: data = 12'h335;
        15'h0BB9: data = 12'h26F;
        15'h0BBA: data = 12'h199;
        15'h0BBB: data = 12'h0B7;
        15'h0BBC: data = 12'h78A;
        15'h0BBD: data = 12'h50D;
        15'h0BBE: data = 12'h58B;
        15'h0BBF: data = 12'h489;
        15'h0BC0: data = 12'h36C;
        15'h0BC1: data = 12'h260;
        15'h0BC2: data = 12'h145;
        15'h0BC3: data = 12'h06F;
        15'h0BC4: data = 12'h6BC;
        15'h0BC5: data = 12'h592;
        15'h0BC6: data = 12'h479;
        15'h0BC7: data = 12'h358;
        15'h0BC8: data = 12'h23D;
        15'h0BC9: data = 12'h128;
        15'h0BCA: data = 12'h027;
        15'h0BCB: data = 12'h6F5;
        15'h0BCC: data = 12'h60C;
        15'h0BCD: data = 12'h52F;
        15'h0BCE: data = 12'h469;
        15'h0BCF: data = 12'h3A0;
        15'h0BD0: data = 12'h2E6;
        15'h0BD1: data = 12'h23D;
        15'h0BD2: data = 12'h1A6;
        15'h0BD3: data = 12'h119;
        15'h0BD4: data = 12'h0BC;
        15'h0BD5: data = 12'h05C;
        15'h0BD6: data = 12'h7A6;
        15'h0BD7: data = 12'h773;
        15'h0BD8: data = 12'h76D;
        15'h0BD9: data = 12'h757;
        15'h0BDA: data = 12'h780;
        15'h0BDB: data = 12'h7A6;
        15'h0BDC: data = 12'h50D;
        15'h0BDD: data = 12'h09C;
        15'h0BDE: data = 12'h10A;
        15'h0BDF: data = 12'h179;
        15'h0BE0: data = 12'h20D;
        15'h0BE1: data = 12'h2A9;
        15'h0BE2: data = 12'h35C;
        15'h0BE3: data = 12'h426;
        15'h0BE4: data = 12'h4F7;
        15'h0BE5: data = 12'h5E1;
        15'h0BE6: data = 12'h6D8;
        15'h0BE7: data = 12'h7CF;
        15'h0BE8: data = 12'h107;
        15'h0BE9: data = 12'h210;
        15'h0BEA: data = 12'h31B;
        15'h0BEB: data = 12'h434;
        15'h0BEC: data = 12'h546;
        15'h0BED: data = 12'h667;
        15'h0BEE: data = 12'h786;
        15'h0BEF: data = 12'h0F7;
        15'h0BF0: data = 12'h216;
        15'h0BF1: data = 12'h33D;
        15'h0BF2: data = 12'h455;
        15'h0BF3: data = 12'h564;
        15'h0BF4: data = 12'h663;
        15'h0BF5: data = 12'h762;
        15'h0BF6: data = 12'h46E;
        15'h0BF7: data = 12'h16A;
        15'h0BF8: data = 12'h23A;
        15'h0BF9: data = 12'h2FD;
        15'h0BFA: data = 12'h3B2;
        15'h0BFB: data = 12'h50D;
        15'h0BFC: data = 12'h4EE;
        15'h0BFD: data = 12'h562;
        15'h0BFE: data = 12'h5D4;
        15'h0BFF: data = 12'h615;
        15'h0C00: data = 12'h659;
        15'h0C01: data = 12'h686;
        15'h0C02: data = 12'h68A;
        15'h0C03: data = 12'h68A;
        15'h0C04: data = 12'h666;
        15'h0C05: data = 12'h632;
        15'h0C06: data = 12'h5EB;
        15'h0C07: data = 12'h59B;
        15'h0C08: data = 12'h534;
        15'h0C09: data = 12'h4B0;
        15'h0C0A: data = 12'h41A;
        15'h0C0B: data = 12'h36C;
        15'h0C0C: data = 12'h2B5;
        15'h0C0D: data = 12'h1DF;
        15'h0C0E: data = 12'h102;
        15'h0C0F: data = 12'h018;
        15'h0C10: data = 12'h6E2;
        15'h0C11: data = 12'h5E5;
        15'h0C12: data = 12'h4DC;
        15'h0C13: data = 12'h3CC;
        15'h0C14: data = 12'h2B4;
        15'h0C15: data = 12'h1A2;
        15'h0C16: data = 12'h086;
        15'h0C17: data = 12'h70D;
        15'h0C18: data = 12'h5F9;
        15'h0C19: data = 12'h4DB;
        15'h0C1A: data = 12'h50D;
        15'h0C1B: data = 12'h29B;
        15'h0C1C: data = 12'h17F;
        15'h0C1D: data = 12'h07F;
        15'h0C1E: data = 12'h745;
        15'h0C1F: data = 12'h65E;
        15'h0C20: data = 12'h573;
        15'h0C21: data = 12'h4A2;
        15'h0C22: data = 12'h3D9;
        15'h0C23: data = 12'h31B;
        15'h0C24: data = 12'h279;
        15'h0C25: data = 12'h1DC;
        15'h0C26: data = 12'h147;
        15'h0C27: data = 12'h0DF;
        15'h0C28: data = 12'h07D;
        15'h0C29: data = 12'h027;
        15'h0C2A: data = 12'h798;
        15'h0C2B: data = 12'h773;
        15'h0C2C: data = 12'h756;
        15'h0C2D: data = 12'h778;
        15'h0C2E: data = 12'h7A0;
        15'h0C2F: data = 12'h7E0;
        15'h0C30: data = 12'h821;
        15'h0C31: data = 12'h0E5;
        15'h0C32: data = 12'h155;
        15'h0C33: data = 12'h1D9;
        15'h0C34: data = 12'h275;
        15'h0C35: data = 12'h321;
        15'h0C36: data = 12'h3E0;
        15'h0C37: data = 12'h4B1;
        15'h0C38: data = 12'h58C;
        15'h0C39: data = 12'h50D;
        15'h0C3A: data = 12'h777;
        15'h0C3B: data = 12'h0C0;
        15'h0C3C: data = 12'h1AF;
        15'h0C3D: data = 12'h2C7;
        15'h0C3E: data = 12'h3D9;
        15'h0C3F: data = 12'h4F4;
        15'h0C40: data = 12'h606;
        15'h0C41: data = 12'h71C;
        15'h0C42: data = 12'h354;
        15'h0C43: data = 12'h1AE;
        15'h0C44: data = 12'h2D3;
        15'h0C45: data = 12'h3F7;
        15'h0C46: data = 12'h50C;
        15'h0C47: data = 12'h616;
        15'h0C48: data = 12'h70E;
        15'h0C49: data = 12'h7FC;
        15'h0C4A: data = 12'h116;
        15'h0C4B: data = 12'h1E9;
        15'h0C4C: data = 12'h2B7;
        15'h0C4D: data = 12'h373;
        15'h0C4E: data = 12'h41D;
        15'h0C4F: data = 12'h4BB;
        15'h0C50: data = 12'h545;
        15'h0C51: data = 12'h5B3;
        15'h0C52: data = 12'h5FC;
        15'h0C53: data = 12'h64F;
        15'h0C54: data = 12'h671;
        15'h0C55: data = 12'h68A;
        15'h0C56: data = 12'h684;
        15'h0C57: data = 12'h664;
        15'h0C58: data = 12'h50D;
        15'h0C59: data = 12'h607;
        15'h0C5A: data = 12'h5BF;
        15'h0C5B: data = 12'h557;
        15'h0C5C: data = 12'h4DD;
        15'h0C5D: data = 12'h453;
        15'h0C5E: data = 12'h3A9;
        15'h0C5F: data = 12'h2F2;
        15'h0C60: data = 12'h22B;
        15'h0C61: data = 12'h14C;
        15'h0C62: data = 12'h067;
        15'h0C63: data = 12'h735;
        15'h0C64: data = 12'h635;
        15'h0C65: data = 12'h530;
        15'h0C66: data = 12'h425;
        15'h0C67: data = 12'h31B;
        15'h0C68: data = 12'h1FF;
        15'h0C69: data = 12'h0E5;
        15'h0C6A: data = 12'h77F;
        15'h0C6B: data = 12'h653;
        15'h0C6C: data = 12'h530;
        15'h0C6D: data = 12'h417;
        15'h0C6E: data = 12'h2F6;
        15'h0C6F: data = 12'h1DC;
        15'h0C70: data = 12'h0D1;
        15'h0C71: data = 12'h7A3;
        15'h0C72: data = 12'h6AB;
        15'h0C73: data = 12'h5C2;
        15'h0C74: data = 12'h4E9;
        15'h0C75: data = 12'h418;
        15'h0C76: data = 12'h357;
        15'h0C77: data = 12'h50D;
        15'h0C78: data = 12'h206;
        15'h0C79: data = 12'h17A;
        15'h0C7A: data = 12'h101;
        15'h0C7B: data = 12'h09A;
        15'h0C7C: data = 12'h03A;
        15'h0C7D: data = 12'h792;
        15'h0C7E: data = 12'h775;
        15'h0C7F: data = 12'h755;
        15'h0C80: data = 12'h777;
        15'h0C81: data = 12'h780;
        15'h0C82: data = 12'h7C3;
        15'h0C83: data = 12'h804;
        15'h0C84: data = 12'h0C2;
        15'h0C85: data = 12'h128;
        15'h0C86: data = 12'h1B3;
        15'h0C87: data = 12'h242;
        15'h0C88: data = 12'h2E6;
        15'h0C89: data = 12'h39F;
        15'h0C8A: data = 12'h469;
        15'h0C8B: data = 12'h53F;
        15'h0C8C: data = 12'h62A;
        15'h0C8D: data = 12'h722;
        15'h0C8E: data = 12'h825;
        15'h0C8F: data = 12'h15C;
        15'h0C90: data = 12'h269;
        15'h0C91: data = 12'h37E;
        15'h0C92: data = 12'h495;
        15'h0C93: data = 12'h5A3;
        15'h0C94: data = 12'h6CB;
        15'h0C95: data = 12'h7E0;
        15'h0C96: data = 12'h50D;
        15'h0C97: data = 12'h277;
        15'h0C98: data = 12'h395;
        15'h0C99: data = 12'h4B4;
        15'h0C9A: data = 12'h5B9;
        15'h0C9B: data = 12'h6C2;
        15'h0C9C: data = 12'h7B1;
        15'h0C9D: data = 12'h0D5;
        15'h0C9E: data = 12'h1AB;
        15'h0C9F: data = 12'h279;
        15'h0CA0: data = 12'h335;
        15'h0CA1: data = 12'h3E9;
        15'h0CA2: data = 12'h490;
        15'h0CA3: data = 12'h519;
        15'h0CA4: data = 12'h58A;
        15'h0CA5: data = 12'h5F4;
        15'h0CA6: data = 12'h638;
        15'h0CA7: data = 12'h670;
        15'h0CA8: data = 12'h68D;
        15'h0CA9: data = 12'h688;
        15'h0CAA: data = 12'h686;
        15'h0CAB: data = 12'h664;
        15'h0CAC: data = 12'h623;
        15'h0CAD: data = 12'h5D3;
        15'h0CAE: data = 12'h56D;
        15'h0CAF: data = 12'h50A;
        15'h0CB0: data = 12'h481;
        15'h0CB1: data = 12'h3E7;
        15'h0CB2: data = 12'h335;
        15'h0CB3: data = 12'h271;
        15'h0CB4: data = 12'h199;
        15'h0CB5: data = 12'h50D;
        15'h0CB6: data = 12'h78A;
        15'h0CB7: data = 12'h692;
        15'h0CB8: data = 12'h589;
        15'h0CB9: data = 12'h488;
        15'h0CBA: data = 12'h36A;
        15'h0CBB: data = 12'h258;
        15'h0CBC: data = 12'h140;
        15'h0CBD: data = 12'h0E7;
        15'h0CBE: data = 12'h6B9;
        15'h0CBF: data = 12'h591;
        15'h0CC0: data = 12'h47B;
        15'h0CC1: data = 12'h35F;
        15'h0CC2: data = 12'h240;
        15'h0CC3: data = 12'h128;
        15'h0CC4: data = 12'h02A;
        15'h0CC5: data = 12'h6F3;
        15'h0CC6: data = 12'h601;
        15'h0CC7: data = 12'h528;
        15'h0CC8: data = 12'h45A;
        15'h0CC9: data = 12'h397;
        15'h0CCA: data = 12'h2E5;
        15'h0CCB: data = 12'h23D;
        15'h0CCC: data = 12'h1A8;
        15'h0CCD: data = 12'h11B;
        15'h0CCE: data = 12'h0BF;
        15'h0CCF: data = 12'h05B;
        15'h0CD0: data = 12'h79D;
        15'h0CD1: data = 12'h770;
        15'h0CD2: data = 12'h767;
        15'h0CD3: data = 12'h74E;
        15'h0CD4: data = 12'h50D;
        15'h0CD5: data = 12'h79F;
        15'h0CD6: data = 12'h7ED;
        15'h0CD7: data = 12'h0AC;
        15'h0CD8: data = 12'h108;
        15'h0CD9: data = 12'h17D;
        15'h0CDA: data = 12'h20F;
        15'h0CDB: data = 12'h2AF;
        15'h0CDC: data = 12'h35E;
        15'h0CDD: data = 12'h420;
        15'h0CDE: data = 12'h4F8;
        15'h0CDF: data = 12'h5DC;
        15'h0CE0: data = 12'h6CE;
        15'h0CE1: data = 12'h7C7;
        15'h0CE2: data = 12'h101;
        15'h0CE3: data = 12'h20E;
        15'h0CE4: data = 12'h31B;
        15'h0CE5: data = 12'h43C;
        15'h0CE6: data = 12'h54B;
        15'h0CE7: data = 12'h66B;
        15'h0CE8: data = 12'h786;
        15'h0CE9: data = 12'h0F4;
        15'h0CEA: data = 12'h20C;
        15'h0CEB: data = 12'h32C;
        15'h0CEC: data = 12'h44E;
        15'h0CED: data = 12'h55D;
        15'h0CEE: data = 12'h669;
        15'h0CEF: data = 12'h763;
        15'h0CF0: data = 12'h574;
        15'h0CF1: data = 12'h16D;
        15'h0CF2: data = 12'h237;
        15'h0CF3: data = 12'h50D;
        15'h0CF4: data = 12'h3AE;
        15'h0CF5: data = 12'h44B;
        15'h0CF6: data = 12'h4E4;
        15'h0CF7: data = 12'h55A;
        15'h0CF8: data = 12'h5D1;
        15'h0CF9: data = 12'h615;
        15'h0CFA: data = 12'h656;
        15'h0CFB: data = 12'h688;
        15'h0CFC: data = 12'h695;
        15'h0CFD: data = 12'h68D;
        15'h0CFE: data = 12'h664;
        15'h0CFF: data = 12'h632;
        15'h0D00: data = 12'h5E0;
        15'h0D01: data = 12'h58F;
        15'h0D02: data = 12'h52E;
        15'h0D03: data = 12'h4A9;
        15'h0D04: data = 12'h413;
        15'h0D05: data = 12'h36A;
        15'h0D06: data = 12'h2B1;
        15'h0D07: data = 12'h1E4;
        15'h0D08: data = 12'h10D;
        15'h0D09: data = 12'h020;
        15'h0D0A: data = 12'h6E5;
        15'h0D0B: data = 12'h5E3;
        15'h0D0C: data = 12'h4D8;
        15'h0D0D: data = 12'h3C5;
        15'h0D0E: data = 12'h2AB;
        15'h0D0F: data = 12'h192;
        15'h0D10: data = 12'h07E;
        15'h0D11: data = 12'h70E;
        15'h0D12: data = 12'h50D;
        15'h0D13: data = 12'h4E2;
        15'h0D14: data = 12'h3BA;
        15'h0D15: data = 12'h2A5;
        15'h0D16: data = 12'h18A;
        15'h0D17: data = 12'h082;
        15'h0D18: data = 12'h745;
        15'h0D19: data = 12'h65C;
        15'h0D1A: data = 12'h569;
        15'h0D1B: data = 12'h499;
        15'h0D1C: data = 12'h3CC;
        15'h0D1D: data = 12'h316;
        15'h0D1E: data = 12'h273;
        15'h0D1F: data = 12'h1D9;
        15'h0D20: data = 12'h147;
        15'h0D21: data = 12'h0E6;
        15'h0D22: data = 12'h088;
        15'h0D23: data = 12'h039;
        15'h0D24: data = 12'h79B;
        15'h0D25: data = 12'h775;
        15'h0D26: data = 12'h755;
        15'h0D27: data = 12'h776;
        15'h0D28: data = 12'h796;
        15'h0D29: data = 12'h7D2;
        15'h0D2A: data = 12'h81D;
        15'h0D2B: data = 12'h0E5;
        15'h0D2C: data = 12'h152;
        15'h0D2D: data = 12'h1DF;
        15'h0D2E: data = 12'h27D;
        15'h0D2F: data = 12'h32E;
        15'h0D30: data = 12'h3E7;
        15'h0D31: data = 12'h50D;
        15'h0D32: data = 12'h584;
        15'h0D33: data = 12'h673;
        15'h0D34: data = 12'h766;
        15'h0D35: data = 12'h0F9;
        15'h0D36: data = 12'h1A8;
        15'h0D37: data = 12'h2CB;
        15'h0D38: data = 12'h3DC;
        15'h0D39: data = 12'h4FC;
        15'h0D3A: data = 12'h611;
        15'h0D3B: data = 12'h72A;
        15'h0D3C: data = 12'h4C0;
        15'h0D3D: data = 12'h1AF;
        15'h0D3E: data = 12'h2CB;
        15'h0D3F: data = 12'h3EC;
        15'h0D40: data = 12'h4FD;
        15'h0D41: data = 12'h60E;
        15'h0D42: data = 12'h710;
        15'h0D43: data = 12'h804;
        15'h0D44: data = 12'h125;
        15'h0D45: data = 12'h1FC;
        15'h0D46: data = 12'h2BB;
        15'h0D47: data = 12'h372;
        15'h0D48: data = 12'h416;
        15'h0D49: data = 12'h4B0;
        15'h0D4A: data = 12'h537;
        15'h0D4B: data = 12'h5A4;
        15'h0D4C: data = 12'h5F1;
        15'h0D4D: data = 12'h653;
        15'h0D4E: data = 12'h677;
        15'h0D4F: data = 12'h698;
        15'h0D50: data = 12'h50D;
        15'h0D51: data = 12'h674;
        15'h0D52: data = 12'h64E;
        15'h0D53: data = 12'h609;
        15'h0D54: data = 12'h5B1;
        15'h0D55: data = 12'h54C;
        15'h0D56: data = 12'h4CC;
        15'h0D57: data = 12'h446;
        15'h0D58: data = 12'h3A4;
        15'h0D59: data = 12'h2F2;
        15'h0D5A: data = 12'h22D;
        15'h0D5B: data = 12'h152;
        15'h0D5C: data = 12'h074;
        15'h0D5D: data = 12'h73E;
        15'h0D5E: data = 12'h641;
        15'h0D5F: data = 12'h53C;
        15'h0D60: data = 12'h422;
        15'h0D61: data = 12'h311;
        15'h0D62: data = 12'h1F1;
        15'h0D63: data = 12'h0D7;
        15'h0D64: data = 12'h771;
        15'h0D65: data = 12'h64B;
        15'h0D66: data = 12'h52F;
        15'h0D67: data = 12'h41F;
        15'h0D68: data = 12'h301;
        15'h0D69: data = 12'h1EE;
        15'h0D6A: data = 12'h0DE;
        15'h0D6B: data = 12'h788;
        15'h0D6C: data = 12'h6AB;
        15'h0D6D: data = 12'h5C0;
        15'h0D6E: data = 12'h4E4;
        15'h0D6F: data = 12'h50D;
        15'h0D70: data = 12'h348;
        15'h0D71: data = 12'h297;
        15'h0D72: data = 12'h1FA;
        15'h0D73: data = 12'h16F;
        15'h0D74: data = 12'h0FF;
        15'h0D75: data = 12'h0A1;
        15'h0D76: data = 12'h046;
        15'h0D77: data = 12'h7A0;
        15'h0D78: data = 12'h780;
        15'h0D79: data = 12'h75D;
        15'h0D7A: data = 12'h775;
        15'h0D7B: data = 12'h772;
        15'h0D7C: data = 12'h7B0;
        15'h0D7D: data = 12'h7F4;
        15'h0D7E: data = 12'h0B9;
        15'h0D7F: data = 12'h121;
        15'h0D80: data = 12'h1B2;
        15'h0D81: data = 12'h24E;
        15'h0D82: data = 12'h2F5;
        15'h0D83: data = 12'h3AD;
        15'h0D84: data = 12'h47A;
        15'h0D85: data = 12'h543;
        15'h0D86: data = 12'h628;
        15'h0D87: data = 12'h713;
        15'h0D88: data = 12'h80F;
        15'h0D89: data = 12'h14A;
        15'h0D8A: data = 12'h25D;
        15'h0D8B: data = 12'h37D;
        15'h0D8C: data = 12'h49C;
        15'h0D8D: data = 12'h5B2;
        15'h0D8E: data = 12'h50D;
        15'h0D8F: data = 12'h7F4;
        15'h0D90: data = 12'h156;
        15'h0D91: data = 12'h274;
        15'h0D92: data = 12'h385;
        15'h0D93: data = 12'h4A2;
        15'h0D94: data = 12'h5A9;
        15'h0D95: data = 12'h6B7;
        15'h0D96: data = 12'h7AF;
        15'h0D97: data = 12'h0E3;
        15'h0D98: data = 12'h1BB;
        15'h0D99: data = 12'h28C;
        15'h0D9A: data = 12'h340;
        15'h0D9B: data = 12'h3F2;
        15'h0D9C: data = 12'h48A;
        15'h0D9D: data = 12'h50B;
        15'h0D9E: data = 12'h57B;
        15'h0D9F: data = 12'h5E3;
        15'h0DA0: data = 12'h628;
        15'h0DA1: data = 12'h66E;
        15'h0DA2: data = 12'h691;
        15'h0DA3: data = 12'h695;
        15'h0DA4: data = 12'h694;
        15'h0DA5: data = 12'h670;
        15'h0DA6: data = 12'h634;
        15'h0DA7: data = 12'h5D9;
        15'h0DA8: data = 12'h567;
        15'h0DA9: data = 12'h4F6;
        15'h0DAA: data = 12'h469;
        15'h0DAB: data = 12'h3D1;
        15'h0DAC: data = 12'h326;
        15'h0DAD: data = 12'h50D;
        15'h0DAE: data = 12'h19A;
        15'h0DAF: data = 12'h0C5;
        15'h0DB0: data = 12'h791;
        15'h0DB1: data = 12'h6A3;
        15'h0DB2: data = 12'h598;
        15'h0DB3: data = 12'h48F;
        15'h0DB4: data = 12'h367;
        15'h0DB5: data = 12'h252;
        15'h0DB6: data = 12'h132;
        15'h0DB7: data = 12'h01E;
        15'h0DB8: data = 12'h6A7;
        15'h0DB9: data = 12'h584;
        15'h0DBA: data = 12'h470;
        15'h0DBB: data = 12'h358;
        15'h0DBC: data = 12'h247;
        15'h0DBD: data = 12'h131;
        15'h0DBE: data = 12'h036;
        15'h0DBF: data = 12'h706;
        15'h0DC0: data = 12'h615;
        15'h0DC1: data = 12'h531;
        15'h0DC2: data = 12'h45E;
        15'h0DC3: data = 12'h38B;
        15'h0DC4: data = 12'h2D0;
        15'h0DC5: data = 12'h229;
        15'h0DC6: data = 12'h199;
        15'h0DC7: data = 12'h110;
        15'h0DC8: data = 12'h0C1;
        15'h0DC9: data = 12'h067;
        15'h0DCA: data = 12'h733;
        15'h0DCB: data = 12'h783;
        15'h0DCC: data = 12'h50D;
        15'h0DCD: data = 12'h75F;
        15'h0DCE: data = 12'h779;
        15'h0DCF: data = 12'h79A;
        15'h0DD0: data = 12'h7DD;
        15'h0DD1: data = 12'h093;
        15'h0DD2: data = 12'h0FC;
        15'h0DD3: data = 12'h174;
        15'h0DD4: data = 12'h20F;
        15'h0DD5: data = 12'h2B3;
        15'h0DD6: data = 12'h371;
        15'h0DD7: data = 12'h435;
        15'h0DD8: data = 12'h508;
        15'h0DD9: data = 12'h5EA;
        15'h0DDA: data = 12'h6D5;
        15'h0DDB: data = 12'h7C7;
        15'h0DDC: data = 12'h0F9;
        15'h0DDD: data = 12'h1FF;
        15'h0DDE: data = 12'h305;
        15'h0DDF: data = 12'h42C;
        15'h0DE0: data = 12'h54B;
        15'h0DE1: data = 12'h677;
        15'h0DE2: data = 12'h79A;
        15'h0DE3: data = 12'h102;
        15'h0DE4: data = 12'h21D;
        15'h0DE5: data = 12'h331;
        15'h0DE6: data = 12'h444;
        15'h0DE7: data = 12'h54F;
        15'h0DE8: data = 12'h657;
        15'h0DE9: data = 12'h755;
        15'h0DEA: data = 12'h1A6;
        15'h0DEB: data = 12'h50D;
        15'h0DEC: data = 12'h243;
        15'h0DED: data = 12'h306;
        15'h0DEE: data = 12'h3BE;
        15'h0DEF: data = 12'h45A;
        15'h0DF0: data = 12'h4F1;
        15'h0DF1: data = 12'h55B;
        15'h0DF2: data = 12'h5C8;
        15'h0DF3: data = 12'h607;
        15'h0DF4: data = 12'h649;
        15'h0DF5: data = 12'h67F;
        15'h0DF6: data = 12'h68E;
        15'h0DF7: data = 12'h692;
        15'h0DF8: data = 12'h675;
        15'h0DF9: data = 12'h642;
        15'h0DFA: data = 12'h5F4;
        15'h0DFB: data = 12'h59F;
        15'h0DFC: data = 12'h537;
        15'h0DFD: data = 12'h4A6;
        15'h0DFE: data = 12'h408;
        15'h0DFF: data = 12'h358;
        15'h0E00: data = 12'h2A3;
        15'h0E01: data = 12'h1D8;
        15'h0E02: data = 12'h108;
        15'h0E03: data = 12'h0A8;
        15'h0E04: data = 12'h6F1;
        15'h0E05: data = 12'h5F4;
        15'h0E06: data = 12'h4E7;
        15'h0E07: data = 12'h3D7;
        15'h0E08: data = 12'h2BB;
        15'h0E09: data = 12'h1A2;
        15'h0E0A: data = 12'h50D;
        15'h0E0B: data = 12'h6FE;
        15'h0E0C: data = 12'h5EA;
        15'h0E0D: data = 12'h4D2;
        15'h0E0E: data = 12'h3AD;
        15'h0E0F: data = 12'h29A;
        15'h0E10: data = 12'h189;
        15'h0E11: data = 12'h08A;
        15'h0E12: data = 12'h750;
        15'h0E13: data = 12'h66F;
        15'h0E14: data = 12'h57C;
        15'h0E15: data = 12'h4A9;
        15'h0E16: data = 12'h3D7;
        15'h0E17: data = 12'h315;
        15'h0E18: data = 12'h25F;
        15'h0E19: data = 12'h1C5;
        15'h0E1A: data = 12'h136;
        15'h0E1B: data = 12'h0D7;
        15'h0E1C: data = 12'h07C;
        15'h0E1D: data = 12'h031;
        15'h0E1E: data = 12'h7A7;
        15'h0E1F: data = 12'h784;
        15'h0E20: data = 12'h763;
        15'h0E21: data = 12'h784;
        15'h0E22: data = 12'h79E;
        15'h0E23: data = 12'h7D9;
        15'h0E24: data = 12'h571;
        15'h0E25: data = 12'h0D7;
        15'h0E26: data = 12'h147;
        15'h0E27: data = 12'h1CF;
        15'h0E28: data = 12'h26A;
        15'h0E29: data = 12'h50D;
        15'h0E2A: data = 12'h3EA;
        15'h0E2B: data = 12'h4BC;
        15'h0E2C: data = 12'h59A;
        15'h0E2D: data = 12'h687;
        15'h0E2E: data = 12'h77B;
        15'h0E2F: data = 12'h0AA;
        15'h0E30: data = 12'h19F;
        15'h0E31: data = 12'h2B8;
        15'h0E32: data = 12'h3CD;
        15'h0E33: data = 12'h4F1;
        15'h0E34: data = 12'h60A;
        15'h0E35: data = 12'h72A;
        15'h0E36: data = 12'h659;
        15'h0E37: data = 12'h1C2;
        15'h0E38: data = 12'h2DF;
        15'h0E39: data = 12'h3F5;
        15'h0E3A: data = 12'h500;
        15'h0E3B: data = 12'h603;
        15'h0E3C: data = 12'h702;
        15'h0E3D: data = 12'h7F4;
        15'h0E3E: data = 12'h11D;
        15'h0E3F: data = 12'h1F5;
        15'h0E40: data = 12'h2C5;
        15'h0E41: data = 12'h380;
        15'h0E42: data = 12'h427;
        15'h0E43: data = 12'h4BF;
        15'h0E44: data = 12'h544;
        15'h0E45: data = 12'h5AB;
        15'h0E46: data = 12'h5F0;
        15'h0E47: data = 12'h643;
        15'h0E48: data = 12'h50D;
        15'h0E49: data = 12'h684;
        15'h0E4A: data = 12'h688;
        15'h0E4B: data = 12'h672;
        15'h0E4C: data = 12'h653;
        15'h0E4D: data = 12'h616;
        15'h0E4E: data = 12'h5C6;
        15'h0E4F: data = 12'h55A;
        15'h0E50: data = 12'h4DA;
        15'h0E51: data = 12'h44C;
        15'h0E52: data = 12'h39F;
        15'h0E53: data = 12'h2E6;
        15'h0E54: data = 12'h21B;
        15'h0E55: data = 12'h141;
        15'h0E56: data = 12'h065;
        15'h0E57: data = 12'h736;
        15'h0E58: data = 12'h641;
        15'h0E59: data = 12'h542;
        15'h0E5A: data = 12'h430;
        15'h0E5B: data = 12'h328;
        15'h0E5C: data = 12'h201;
        15'h0E5D: data = 12'h0E3;
        15'h0E5E: data = 12'h774;
        15'h0E5F: data = 12'h649;
        15'h0E60: data = 12'h51F;
        15'h0E61: data = 12'h408;
        15'h0E62: data = 12'h2EC;
        15'h0E63: data = 12'h1D6;
        15'h0E64: data = 12'h0D5;
        15'h0E65: data = 12'h7AB;
        15'h0E66: data = 12'h6B5;
        15'h0E67: data = 12'h50D;
        15'h0E68: data = 12'h4F3;
        15'h0E69: data = 12'h41B;
        15'h0E6A: data = 12'h356;
        15'h0E6B: data = 12'h2A0;
        15'h0E6C: data = 12'h1FA;
        15'h0E6D: data = 12'h16D;
        15'h0E6E: data = 12'h0F7;
        15'h0E6F: data = 12'h095;
        15'h0E70: data = 12'h038;
        15'h0E71: data = 12'h798;
        15'h0E72: data = 12'h77C;
        15'h0E73: data = 12'h760;
        15'h0E74: data = 12'h783;
        15'h0E75: data = 12'h789;
        15'h0E76: data = 12'h7C6;
        15'h0E77: data = 12'h803;
        15'h0E78: data = 12'h0C1;
        15'h0E79: data = 12'h11E;
        15'h0E7A: data = 12'h1A7;
        15'h0E7B: data = 12'h23B;
        15'h0E7C: data = 12'h2E7;
        15'h0E7D: data = 12'h3A1;
        15'h0E7E: data = 12'h477;
        15'h0E7F: data = 12'h54A;
        15'h0E80: data = 12'h63B;
        15'h0E81: data = 12'h726;
        15'h0E82: data = 12'h823;
        15'h0E83: data = 12'h155;
        15'h0E84: data = 12'h261;
        15'h0E85: data = 12'h375;
        15'h0E86: data = 12'h50D;
        15'h0E87: data = 12'h5A2;
        15'h0E88: data = 12'h6CD;
        15'h0E89: data = 12'h7EA;
        15'h0E8A: data = 12'h159;
        15'h0E8B: data = 12'h285;
        15'h0E8C: data = 12'h39B;
        15'h0E8D: data = 12'h4B1;
        15'h0E8E: data = 12'h5B3;
        15'h0E8F: data = 12'h6B8;
        15'h0E90: data = 12'h7A4;
        15'h0E91: data = 12'h0D2;
        15'h0E92: data = 12'h1AC;
        15'h0E93: data = 12'h27C;
        15'h0E94: data = 12'h336;
        15'h0E95: data = 12'h3F5;
        15'h0E96: data = 12'h498;
        15'h0E97: data = 12'h520;
        15'h0E98: data = 12'h58A;
        15'h0E99: data = 12'h5F4;
        15'h0E9A: data = 12'h637;
        15'h0E9B: data = 12'h671;
        15'h0E9C: data = 12'h686;
        15'h0E9D: data = 12'h688;
        15'h0E9E: data = 12'h683;
        15'h0E9F: data = 12'h665;
        15'h0EA0: data = 12'h62A;
        15'h0EA1: data = 12'h5DC;
        15'h0EA2: data = 12'h576;
        15'h0EA3: data = 12'h509;
        15'h0EA4: data = 12'h484;
        15'h0EA5: data = 12'h50D;
        15'h0EA6: data = 12'h331;
        15'h0EA7: data = 12'h26A;
        15'h0EA8: data = 12'h192;
        15'h0EA9: data = 12'h0B3;
        15'h0EAA: data = 12'h789;
        15'h0EAB: data = 12'h68E;
        15'h0EAC: data = 12'h58B;
        15'h0EAD: data = 12'h487;
        15'h0EAE: data = 12'h36E;
        15'h0EAF: data = 12'h25E;
        15'h0EB0: data = 12'h143;
        15'h0EB1: data = 12'h022;
        15'h0EB2: data = 12'h6C4;
        15'h0EB3: data = 12'h58D;
        15'h0EB4: data = 12'h474;
        15'h0EB5: data = 12'h352;
        15'h0EB6: data = 12'h238;
        15'h0EB7: data = 12'h121;
        15'h0EB8: data = 12'h028;
        15'h0EB9: data = 12'h6F7;
        15'h0EBA: data = 12'h609;
        15'h0EBB: data = 12'h52B;
        15'h0EBC: data = 12'h462;
        15'h0EBD: data = 12'h39C;
        15'h0EBE: data = 12'h2E1;
        15'h0EBF: data = 12'h23B;
        15'h0EC0: data = 12'h1A4;
        15'h0EC1: data = 12'h116;
        15'h0EC2: data = 12'h0B9;
        15'h0EC3: data = 12'h059;
        15'h0EC4: data = 12'h50D;
        15'h0EC5: data = 12'h774;
        15'h0EC6: data = 12'h769;
        15'h0EC7: data = 12'h759;
        15'h0EC8: data = 12'h77E;
        15'h0EC9: data = 12'h7A6;
        15'h0ECA: data = 12'h7E8;
        15'h0ECB: data = 12'h09C;
        15'h0ECC: data = 12'h10B;
        15'h0ECD: data = 12'h17F;
        15'h0ECE: data = 12'h20D;
        15'h0ECF: data = 12'h2AB;
        15'h0ED0: data = 12'h360;
        15'h0ED1: data = 12'h424;
        15'h0ED2: data = 12'h4F9;
        15'h0ED3: data = 12'h5DF;
        15'h0ED4: data = 12'h6D4;
        15'h0ED5: data = 12'h7CF;
        15'h0ED6: data = 12'h108;
        15'h0ED7: data = 12'h210;
        15'h0ED8: data = 12'h31D;
        15'h0ED9: data = 12'h435;
        15'h0EDA: data = 12'h547;
        15'h0EDB: data = 12'h668;
        15'h0EDC: data = 12'h788;
        15'h0EDD: data = 12'h0F7;
        15'h0EDE: data = 12'h212;
        15'h0EDF: data = 12'h339;
        15'h0EE0: data = 12'h454;
        15'h0EE1: data = 12'h561;
        15'h0EE2: data = 12'h668;
        15'h0EE3: data = 12'h50D;
        15'h0EE4: data = 12'h4BB;
        15'h0EE5: data = 12'h16D;
        15'h0EE6: data = 12'h238;
        15'h0EE7: data = 12'h2F8;
        15'h0EE8: data = 12'h3AF;
        15'h0EE9: data = 12'h454;
        15'h0EEA: data = 12'h4EA;
        15'h0EEB: data = 12'h565;
        15'h0EEC: data = 12'h5D7;
        15'h0EED: data = 12'h619;
        15'h0EEE: data = 12'h657;
        15'h0EEF: data = 12'h685;
        15'h0EF0: data = 12'h68E;
        15'h0EF1: data = 12'h68C;
        15'h0EF2: data = 12'h667;
        15'h0EF3: data = 12'h634;
        15'h0EF4: data = 12'h5E7;
        15'h0EF5: data = 12'h596;
        15'h0EF6: data = 12'h532;
        15'h0EF7: data = 12'h4B0;
        15'h0EF8: data = 12'h419;
        15'h0EF9: data = 12'h36F;
        15'h0EFA: data = 12'h2B6;
        15'h0EFB: data = 12'h1E7;
        15'h0EFC: data = 12'h10B;
        15'h0EFD: data = 12'h01D;
        15'h0EFE: data = 12'h6E8;
        15'h0EFF: data = 12'h5E8;
        15'h0F00: data = 12'h4DA;
        15'h0F01: data = 12'h3C7;
        15'h0F02: data = 12'h50D;
        15'h0F03: data = 12'h19B;
        15'h0F04: data = 12'h084;
        15'h0F05: data = 12'h710;
        15'h0F06: data = 12'h5FA;
        15'h0F07: data = 12'h4E5;
        15'h0F08: data = 12'h3BB;
        15'h0F09: data = 12'h2A1;
        15'h0F0A: data = 12'h186;
        15'h0F0B: data = 12'h080;
        15'h0F0C: data = 12'h746;
        15'h0F0D: data = 12'h660;
        15'h0F0E: data = 12'h56C;
        15'h0F0F: data = 12'h49D;
        15'h0F10: data = 12'h3D9;
        15'h0F11: data = 12'h31E;
        15'h0F12: data = 12'h274;
        15'h0F13: data = 12'h1DC;
        15'h0F14: data = 12'h149;
        15'h0F15: data = 12'h0E6;
        15'h0F16: data = 12'h081;
        15'h0F17: data = 12'h02A;
        15'h0F18: data = 12'h796;
        15'h0F19: data = 12'h771;
        15'h0F1A: data = 12'h752;
        15'h0F1B: data = 12'h775;
        15'h0F1C: data = 12'h7A0;
        15'h0F1D: data = 12'h7DF;
        15'h0F1E: data = 12'h823;
        15'h0F1F: data = 12'h0E9;
        15'h0F20: data = 12'h157;
        15'h0F21: data = 12'h50D;
        15'h0F22: data = 12'h276;
        15'h0F23: data = 12'h327;
        15'h0F24: data = 12'h3E1;
        15'h0F25: data = 12'h4B1;
        15'h0F26: data = 12'h588;
        15'h0F27: data = 12'h681;
        15'h0F28: data = 12'h771;
        15'h0F29: data = 12'h0C9;
        15'h0F2A: data = 12'h1AA;
        15'h0F2B: data = 12'h2C9;
        15'h0F2C: data = 12'h3D9;
        15'h0F2D: data = 12'h4F9;
        15'h0F2E: data = 12'h60E;
        15'h0F2F: data = 12'h721;
        15'h0F30: data = 12'h37E;
        15'h0F31: data = 12'h1AD;
        15'h0F32: data = 12'h2D3;
        15'h0F33: data = 12'h3F4;
        15'h0F34: data = 12'h50A;
        15'h0F35: data = 12'h613;
        15'h0F36: data = 12'h714;
        15'h0F37: data = 12'h803;
        15'h0F38: data = 12'h124;
        15'h0F39: data = 12'h1F3;
        15'h0F3A: data = 12'h2B9;
        15'h0F3B: data = 12'h36E;
        15'h0F3C: data = 12'h417;
        15'h0F3D: data = 12'h4B0;
        15'h0F3E: data = 12'h53E;
        15'h0F3F: data = 12'h5B1;
        15'h0F40: data = 12'h50D;
        15'h0F41: data = 12'h656;
        15'h0F42: data = 12'h67B;
        15'h0F43: data = 12'h691;
        15'h0F44: data = 12'h68E;
        15'h0F45: data = 12'h669;
        15'h0F46: data = 12'h645;
        15'h0F47: data = 12'h607;
        15'h0F48: data = 12'h5B7;
        15'h0F49: data = 12'h555;
        15'h0F4A: data = 12'h4D9;
        15'h0F4B: data = 12'h451;
        15'h0F4C: data = 12'h3A8;
        15'h0F4D: data = 12'h2F8;
        15'h0F4E: data = 12'h229;
        15'h0F4F: data = 12'h152;
        15'h0F50: data = 12'h072;
        15'h0F51: data = 12'h73C;
        15'h0F52: data = 12'h63C;
        15'h0F53: data = 12'h533;
        15'h0F54: data = 12'h422;
        15'h0F55: data = 12'h312;
        15'h0F56: data = 12'h1F3;
        15'h0F57: data = 12'h0E2;
        15'h0F58: data = 12'h77B;
        15'h0F59: data = 12'h656;
        15'h0F5A: data = 12'h539;
        15'h0F5B: data = 12'h41D;
        15'h0F5C: data = 12'h2FD;
        15'h0F5D: data = 12'h1E0;
        15'h0F5E: data = 12'h0D4;
        15'h0F5F: data = 12'h50D;
        15'h0F60: data = 12'h6A4;
        15'h0F61: data = 12'h5BD;
        15'h0F62: data = 12'h4E5;
        15'h0F63: data = 12'h413;
        15'h0F64: data = 12'h352;
        15'h0F65: data = 12'h2A5;
        15'h0F66: data = 12'h203;
        15'h0F67: data = 12'h17C;
        15'h0F68: data = 12'h109;
        15'h0F69: data = 12'h0A4;
        15'h0F6A: data = 12'h03E;
        15'h0F6B: data = 12'h794;
        15'h0F6C: data = 12'h775;
        15'h0F6D: data = 12'h753;
        15'h0F6E: data = 12'h776;
        15'h0F6F: data = 12'h779;
        15'h0F70: data = 12'h7BA;
        15'h0F71: data = 12'h802;
        15'h0F72: data = 12'h0C8;
        15'h0F73: data = 12'h12C;
        15'h0F74: data = 12'h1B7;
        15'h0F75: data = 12'h24E;
        15'h0F76: data = 12'h2EE;
        15'h0F77: data = 12'h3A4;
        15'h0F78: data = 12'h46D;
        15'h0F79: data = 12'h53F;
        15'h0F7A: data = 12'h62B;
        15'h0F7B: data = 12'h719;
        15'h0F7C: data = 12'h821;
        15'h0F7D: data = 12'h155;
        15'h0F7E: data = 12'h50D;
        15'h0F7F: data = 12'h384;
        15'h0F80: data = 12'h49F;
        15'h0F81: data = 12'h5B1;
        15'h0F82: data = 12'h6D5;
        15'h0F83: data = 12'h7E8;
        15'h0F84: data = 12'h150;
        15'h0F85: data = 12'h271;
        15'h0F86: data = 12'h391;
        15'h0F87: data = 12'h4AC;
        15'h0F88: data = 12'h5BA;
        15'h0F89: data = 12'h6C6;
        15'h0F8A: data = 12'h7B3;
        15'h0F8B: data = 12'h0DE;
        15'h0F8C: data = 12'h1B9;
        15'h0F8D: data = 12'h280;
        15'h0F8E: data = 12'h330;
        15'h0F8F: data = 12'h3E7;
        15'h0F90: data = 12'h48A;
        15'h0F91: data = 12'h512;
        15'h0F92: data = 12'h586;
        15'h0F93: data = 12'h5F6;
        15'h0F94: data = 12'h63D;
        15'h0F95: data = 12'h67C;
        15'h0F96: data = 12'h692;
        15'h0F97: data = 12'h695;
        15'h0F98: data = 12'h68E;
        15'h0F99: data = 12'h666;
        15'h0F9A: data = 12'h62B;
        15'h0F9B: data = 12'h5D3;
        15'h0F9C: data = 12'h567;
        15'h0F9D: data = 12'h50D;
        15'h0F9E: data = 12'h47A;
        15'h0F9F: data = 12'h3E7;
        15'h0FA0: data = 12'h33A;
        15'h0FA1: data = 12'h276;
        15'h0FA2: data = 12'h19C;
        15'h0FA3: data = 12'h0C3;
        15'h0FA4: data = 12'h78D;
        15'h0FA5: data = 12'h694;
        15'h0FA6: data = 12'h589;
        15'h0FA7: data = 12'h481;
        15'h0FA8: data = 12'h368;
        15'h0FA9: data = 12'h24D;
        15'h0FAA: data = 12'h139;
        15'h0FAB: data = 12'h100;
        15'h0FAC: data = 12'h6B9;
        15'h0FAD: data = 12'h594;
        15'h0FAE: data = 12'h47F;
        15'h0FAF: data = 12'h35F;
        15'h0FB0: data = 12'h248;
        15'h0FB1: data = 12'h12E;
        15'h0FB2: data = 12'h02B;
        15'h0FB3: data = 12'h6F7;
        15'h0FB4: data = 12'h607;
        15'h0FB5: data = 12'h526;
        15'h0FB6: data = 12'h456;
        15'h0FB7: data = 12'h38F;
        15'h0FB8: data = 12'h2DB;
        15'h0FB9: data = 12'h23E;
        15'h0FBA: data = 12'h1AA;
        15'h0FBB: data = 12'h11F;
        15'h0FBC: data = 12'h50D;
        15'h0FBD: data = 12'h065;
        15'h0FBE: data = 12'h78E;
        15'h0FBF: data = 12'h775;
        15'h0FC0: data = 12'h76C;
        15'h0FC1: data = 12'h753;
        15'h0FC2: data = 12'h775;
        15'h0FC3: data = 12'h79C;
        15'h0FC4: data = 12'h7E9;
        15'h0FC5: data = 12'h0D3;
        15'h0FC6: data = 12'h108;
        15'h0FC7: data = 12'h180;
        15'h0FC8: data = 12'h214;
        15'h0FC9: data = 12'h2B5;
        15'h0FCA: data = 12'h36A;
        15'h0FCB: data = 12'h42D;
        15'h0FCC: data = 12'h4FA;
        15'h0FCD: data = 12'h5DA;
        15'h0FCE: data = 12'h6CB;
        15'h0FCF: data = 12'h7C5;
        15'h0FD0: data = 12'h0FD;
        15'h0FD1: data = 12'h211;
        15'h0FD2: data = 12'h31A;
        15'h0FD3: data = 12'h43A;
        15'h0FD4: data = 12'h54D;
        15'h0FD5: data = 12'h66D;
        15'h0FD6: data = 12'h787;
        15'h0FD7: data = 12'h0F5;
        15'h0FD8: data = 12'h20A;
        15'h0FD9: data = 12'h330;
        15'h0FDA: data = 12'h44E;
        15'h0FDB: data = 12'h50D;
        15'h0FDC: data = 12'h665;
        15'h0FDD: data = 12'h760;
        15'h0FDE: data = 12'h5A2;
        15'h0FDF: data = 12'h170;
        15'h0FE0: data = 12'h23E;
        15'h0FE1: data = 12'h2FA;
        15'h0FE2: data = 12'h3B0;
        15'h0FE3: data = 12'h452;
        15'h0FE4: data = 12'h4E6;
        15'h0FE5: data = 12'h558;
        15'h0FE6: data = 12'h5CF;
        15'h0FE7: data = 12'h613;
        15'h0FE8: data = 12'h653;
        15'h0FE9: data = 12'h68B;
        15'h0FEA: data = 12'h695;
        15'h0FEB: data = 12'h692;
        15'h0FEC: data = 12'h670;
        15'h0FED: data = 12'h632;
        15'h0FEE: data = 12'h5E6;
        15'h0FEF: data = 12'h58D;
        15'h0FF0: data = 12'h527;
        15'h0FF1: data = 12'h4A2;
        15'h0FF2: data = 12'h40C;
        15'h0FF3: data = 12'h369;
        15'h0FF4: data = 12'h2B3;
        15'h0FF5: data = 12'h1E5;
        15'h0FF6: data = 12'h10A;
        15'h0FF7: data = 12'h026;
        15'h0FF8: data = 12'h6F0;
        15'h0FF9: data = 12'h5E2;
        15'h0FFA: data = 12'h50D;
        15'h0FFB: data = 12'h3C2;
        15'h0FFC: data = 12'h2A9;
        15'h0FFD: data = 12'h191;
        15'h0FFE: data = 12'h079;
        15'h0FFF: data = 12'h704;
        15'h1000: data = 12'h5F2;
        15'h1001: data = 12'h4DD;
        15'h1002: data = 12'h3B7;
        15'h1003: data = 12'h2A4;
        15'h1004: data = 12'h18D;
        15'h1005: data = 12'h089;
        15'h1006: data = 12'h74A;
        15'h1007: data = 12'h65C;
        15'h1008: data = 12'h56A;
        15'h1009: data = 12'h491;
        15'h100A: data = 12'h3C7;
        15'h100B: data = 12'h30D;
        15'h100C: data = 12'h26D;
        15'h100D: data = 12'h1D7;
        15'h100E: data = 12'h14B;
        15'h100F: data = 12'h0E7;
        15'h1010: data = 12'h088;
        15'h1011: data = 12'h034;
        15'h1012: data = 12'h79F;
        15'h1013: data = 12'h776;
        15'h1014: data = 12'h754;
        15'h1015: data = 12'h76D;
        15'h1016: data = 12'h790;
        15'h1017: data = 12'h7D0;
        15'h1018: data = 12'h81B;
        15'h1019: data = 12'h50D;
        15'h101A: data = 12'h152;
        15'h101B: data = 12'h1DD;
        15'h101C: data = 12'h279;
        15'h101D: data = 12'h332;
        15'h101E: data = 12'h3EF;
        15'h101F: data = 12'h4B9;
        15'h1020: data = 12'h58B;
        15'h1021: data = 12'h67C;
        15'h1022: data = 12'h767;
        15'h1023: data = 12'h100;
        15'h1024: data = 12'h1A1;
        15'h1025: data = 12'h2C5;
        15'h1026: data = 12'h3DE;
        15'h1027: data = 12'h500;
        15'h1028: data = 12'h619;
        15'h1029: data = 12'h733;
        15'h102A: data = 12'h4F0;
        15'h102B: data = 12'h1AE;
        15'h102C: data = 12'h2CD;
        15'h102D: data = 12'h3E8;
        15'h102E: data = 12'h500;
        15'h102F: data = 12'h60A;
        15'h1030: data = 12'h711;
        15'h1031: data = 12'h804;
        15'h1032: data = 12'h129;
        15'h1033: data = 12'h1FE;
        15'h1034: data = 12'h2C9;
        15'h1035: data = 12'h379;
        15'h1036: data = 12'h41F;
        15'h1037: data = 12'h4A7;
        15'h1038: data = 12'h50D;
        15'h1039: data = 12'h5A7;
        15'h103A: data = 12'h5F3;
        15'h103B: data = 12'h652;
        15'h103C: data = 12'h67A;
        15'h103D: data = 12'h696;
        15'h103E: data = 12'h69A;
        15'h103F: data = 12'h675;
        15'h1040: data = 12'h652;
        15'h1041: data = 12'h60A;
        15'h1042: data = 12'h5B0;
        15'h1043: data = 12'h549;
        15'h1044: data = 12'h4CA;
        15'h1045: data = 12'h441;
        15'h1046: data = 12'h39D;
        15'h1047: data = 12'h2F0;
        15'h1048: data = 12'h226;
        15'h1049: data = 12'h156;
        15'h104A: data = 12'h074;
        15'h104B: data = 12'h743;
        15'h104C: data = 12'h644;
        15'h104D: data = 12'h53A;
        15'h104E: data = 12'h427;
        15'h104F: data = 12'h312;
        15'h1050: data = 12'h1F2;
        15'h1051: data = 12'h0D3;
        15'h1052: data = 12'h769;
        15'h1053: data = 12'h644;
        15'h1054: data = 12'h52C;
        15'h1055: data = 12'h41C;
        15'h1056: data = 12'h2FE;
        15'h1057: data = 12'h50D;
        15'h1058: data = 12'h0DE;
        15'h1059: data = 12'h78A;
        15'h105A: data = 12'h6AA;
        15'h105B: data = 12'h5BF;
        15'h105C: data = 12'h4E0;
        15'h105D: data = 12'h40B;
        15'h105E: data = 12'h347;
        15'h105F: data = 12'h29A;
        15'h1060: data = 12'h1F7;
        15'h1061: data = 12'h174;
        15'h1062: data = 12'h103;
        15'h1063: data = 12'h0A5;
        15'h1064: data = 12'h048;
        15'h1065: data = 12'h7A3;
        15'h1066: data = 12'h77F;
        15'h1067: data = 12'h75C;
        15'h1068: data = 12'h775;
        15'h1069: data = 12'h777;
        15'h106A: data = 12'h7B0;
        15'h106B: data = 12'h7F6;
        15'h106C: data = 12'h0B7;
        15'h106D: data = 12'h122;
        15'h106E: data = 12'h1B5;
        15'h106F: data = 12'h24E;
        15'h1070: data = 12'h2F9;
        15'h1071: data = 12'h3B3;
        15'h1072: data = 12'h47D;
        15'h1073: data = 12'h546;
        15'h1074: data = 12'h62C;
        15'h1075: data = 12'h717;
        15'h1076: data = 12'h50D;
        15'h1077: data = 12'h14D;
        15'h1078: data = 12'h263;
        15'h1079: data = 12'h381;
        15'h107A: data = 12'h49C;
        15'h107B: data = 12'h5B4;
        15'h107C: data = 12'h6DC;
        15'h107D: data = 12'h7EF;
        15'h107E: data = 12'h154;
        15'h107F: data = 12'h274;
        15'h1080: data = 12'h38A;
        15'h1081: data = 12'h4A1;
        15'h1082: data = 12'h5AC;
        15'h1083: data = 12'h6BD;
        15'h1084: data = 12'h7B5;
        15'h1085: data = 12'h0DF;
        15'h1086: data = 12'h1B9;
        15'h1087: data = 12'h28C;
        15'h1088: data = 12'h33D;
        15'h1089: data = 12'h3EB;
        15'h108A: data = 12'h487;
        15'h108B: data = 12'h507;
        15'h108C: data = 12'h581;
        15'h108D: data = 12'h5E5;
        15'h108E: data = 12'h632;
        15'h108F: data = 12'h672;
        15'h1090: data = 12'h692;
        15'h1091: data = 12'h697;
        15'h1092: data = 12'h695;
        15'h1093: data = 12'h669;
        15'h1094: data = 12'h632;
        15'h1095: data = 12'h50D;
        15'h1096: data = 12'h567;
        15'h1097: data = 12'h4FB;
        15'h1098: data = 12'h46E;
        15'h1099: data = 12'h3D9;
        15'h109A: data = 12'h331;
        15'h109B: data = 12'h271;
        15'h109C: data = 12'h1A3;
        15'h109D: data = 12'h0C3;
        15'h109E: data = 12'h793;
        15'h109F: data = 12'h69A;
        15'h10A0: data = 12'h591;
        15'h10A1: data = 12'h486;
        15'h10A2: data = 12'h367;
        15'h10A3: data = 12'h24A;
        15'h10A4: data = 12'h137;
        15'h10A5: data = 12'h073;
        15'h10A6: data = 12'h6AD;
        15'h10A7: data = 12'h58A;
        15'h10A8: data = 12'h478;
        15'h10A9: data = 12'h35E;
        15'h10AA: data = 12'h248;
        15'h10AB: data = 12'h131;
        15'h10AC: data = 12'h034;
        15'h10AD: data = 12'h6FF;
        15'h10AE: data = 12'h60D;
        15'h10AF: data = 12'h520;
        15'h10B0: data = 12'h454;
        15'h10B1: data = 12'h389;
        15'h10B2: data = 12'h2D1;
        15'h10B3: data = 12'h231;
        15'h10B4: data = 12'h50D;
        15'h10B5: data = 12'h11E;
        15'h10B6: data = 12'h0C5;
        15'h10B7: data = 12'h066;
        15'h10B8: data = 12'h773;
        15'h10B9: data = 12'h77D;
        15'h10BA: data = 12'h76F;
        15'h10BB: data = 12'h757;
        15'h10BC: data = 12'h774;
        15'h10BD: data = 12'h79A;
        15'h10BE: data = 12'h7DE;
        15'h10BF: data = 12'h09B;
        15'h10C0: data = 12'h106;
        15'h10C1: data = 12'h17F;
        15'h10C2: data = 12'h215;
        15'h10C3: data = 12'h2BA;
        15'h10C4: data = 12'h36F;
        15'h10C5: data = 12'h432;
        15'h10C6: data = 12'h4FE;
        15'h10C7: data = 12'h5DE;
        15'h10C8: data = 12'h6CA;
        15'h10C9: data = 12'h7C1;
        15'h10CA: data = 12'h0F8;
        15'h10CB: data = 12'h205;
        15'h10CC: data = 12'h31C;
        15'h10CD: data = 12'h43D;
        15'h10CE: data = 12'h551;
        15'h10CF: data = 12'h676;
        15'h10D0: data = 12'h799;
        15'h10D1: data = 12'h0FD;
        15'h10D2: data = 12'h210;
        15'h10D3: data = 12'h50D;
        15'h10D4: data = 12'h442;
        15'h10D5: data = 12'h552;
        15'h10D6: data = 12'h65C;
        15'h10D7: data = 12'h75C;
        15'h10D8: data = 12'h3A5;
        15'h10D9: data = 12'h174;
        15'h10DA: data = 12'h245;
        15'h10DB: data = 12'h308;
        15'h10DC: data = 12'h3B8;
        15'h10DD: data = 12'h455;
        15'h10DE: data = 12'h4E2;
        15'h10DF: data = 12'h555;
        15'h10E0: data = 12'h5C3;
        15'h10E1: data = 12'h60C;
        15'h10E2: data = 12'h657;
        15'h10E3: data = 12'h68C;
        15'h10E4: data = 12'h69A;
        15'h10E5: data = 12'h696;
        15'h10E6: data = 12'h675;
        15'h10E7: data = 12'h63C;
        15'h10E8: data = 12'h5EB;
        15'h10E9: data = 12'h58F;
        15'h10EA: data = 12'h527;
        15'h10EB: data = 12'h49D;
        15'h10EC: data = 12'h407;
        15'h10ED: data = 12'h35C;
        15'h10EE: data = 12'h2AB;
        15'h10EF: data = 12'h1E3;
        15'h10F0: data = 12'h10B;
        15'h10F1: data = 12'h029;
        15'h10F2: data = 12'h50D;
        15'h10F3: data = 12'h5ED;
        15'h10F4: data = 12'h4DB;
        15'h10F5: data = 12'h3C5;
        15'h10F6: data = 12'h2A9;
        15'h10F7: data = 12'h18F;
        15'h10F8: data = 12'h06E;
        15'h10F9: data = 12'h6F9;
        15'h10FA: data = 12'h5E3;
        15'h10FB: data = 12'h4D1;
        15'h10FC: data = 12'h3B3;
        15'h10FD: data = 12'h2A5;
        15'h10FE: data = 12'h190;
        15'h10FF: data = 12'h08C;
        15'h1100: data = 12'h74E;
        15'h1101: data = 12'h669;
        15'h1102: data = 12'h570;
        15'h1103: data = 12'h499;
        15'h1104: data = 12'h3C6;
        15'h1105: data = 12'h30A;
        15'h1106: data = 12'h260;
        15'h1107: data = 12'h1CB;
        15'h1108: data = 12'h13B;
        15'h1109: data = 12'h0E3;
        15'h110A: data = 12'h086;
        15'h110B: data = 12'h037;
        15'h110C: data = 12'h7A8;
        15'h110D: data = 12'h782;
        15'h110E: data = 12'h75F;
        15'h110F: data = 12'h777;
        15'h1110: data = 12'h793;
        15'h1111: data = 12'h50D;
        15'h1112: data = 12'h38F;
        15'h1113: data = 12'h0D8;
        15'h1114: data = 12'h14C;
        15'h1115: data = 12'h1D8;
        15'h1116: data = 12'h27C;
        15'h1117: data = 12'h331;
        15'h1118: data = 12'h3EF;
        15'h1119: data = 12'h4BE;
        15'h111A: data = 12'h594;
        15'h111B: data = 12'h67E;
        15'h111C: data = 12'h76D;
        15'h111D: data = 12'h12B;
        15'h111E: data = 12'h19F;
        15'h111F: data = 12'h2BF;
        15'h1120: data = 12'h3D7;
        15'h1121: data = 12'h4FA;
        15'h1122: data = 12'h613;
        15'h1123: data = 12'h72F;
        15'h1124: data = 12'h57B;
        15'h1125: data = 12'h1C1;
        15'h1126: data = 12'h2D6;
        15'h1127: data = 12'h3EE;
        15'h1128: data = 12'h4FB;
        15'h1129: data = 12'h5FF;
        15'h112A: data = 12'h702;
        15'h112B: data = 12'h7FA;
        15'h112C: data = 12'h125;
        15'h112D: data = 12'h1FC;
        15'h112E: data = 12'h2C9;
        15'h112F: data = 12'h380;
        15'h1130: data = 12'h50D;
        15'h1131: data = 12'h4B2;
        15'h1132: data = 12'h534;
        15'h1133: data = 12'h599;
        15'h1134: data = 12'h5EA;
        15'h1135: data = 12'h642;
        15'h1136: data = 12'h66A;
        15'h1137: data = 12'h690;
        15'h1138: data = 12'h693;
        15'h1139: data = 12'h677;
        15'h113A: data = 12'h655;
        15'h113B: data = 12'h60E;
        15'h113C: data = 12'h5B8;
        15'h113D: data = 12'h550;
        15'h113E: data = 12'h4CB;
        15'h113F: data = 12'h43D;
        15'h1140: data = 12'h396;
        15'h1141: data = 12'h2E6;
        15'h1142: data = 12'h220;
        15'h1143: data = 12'h14D;
        15'h1144: data = 12'h075;
        15'h1145: data = 12'h743;
        15'h1146: data = 12'h645;
        15'h1147: data = 12'h544;
        15'h1148: data = 12'h428;
        15'h1149: data = 12'h318;
        15'h114A: data = 12'h1F5;
        15'h114B: data = 12'h0D1;
        15'h114C: data = 12'h76C;
        15'h114D: data = 12'h63D;
        15'h114E: data = 12'h520;
        15'h114F: data = 12'h50D;
        15'h1150: data = 12'h2F8;
        15'h1151: data = 12'h1E4;
        15'h1152: data = 12'h0DF;
        15'h1153: data = 12'h786;
        15'h1154: data = 12'h6B6;
        15'h1155: data = 12'h5C7;
        15'h1156: data = 12'h4EF;
        15'h1157: data = 12'h412;
        15'h1158: data = 12'h347;
        15'h1159: data = 12'h28E;
        15'h115A: data = 12'h1ED;
        15'h115B: data = 12'h166;
        15'h115C: data = 12'h0F6;
        15'h115D: data = 12'h09A;
        15'h115E: data = 12'h042;
        15'h115F: data = 12'h7A5;
        15'h1160: data = 12'h786;
        15'h1161: data = 12'h764;
        15'h1162: data = 12'h77D;
        15'h1163: data = 12'h779;
        15'h1164: data = 12'h7B9;
        15'h1165: data = 12'h7F1;
        15'h1166: data = 12'h0B4;
        15'h1167: data = 12'h116;
        15'h1168: data = 12'h1A7;
        15'h1169: data = 12'h246;
        15'h116A: data = 12'h2F2;
        15'h116B: data = 12'h3AF;
        15'h116C: data = 12'h47B;
        15'h116D: data = 12'h54A;
        15'h116E: data = 12'h50D;
        15'h116F: data = 12'h71B;
        15'h1170: data = 12'h814;
        15'h1171: data = 12'h146;
        15'h1172: data = 12'h255;
        15'h1173: data = 12'h372;
        15'h1174: data = 12'h493;
        15'h1175: data = 12'h5AB;
        15'h1176: data = 12'h6DB;
        15'h1177: data = 12'h7F2;
        15'h1178: data = 12'h15E;
        15'h1179: data = 12'h27D;
        15'h117A: data = 12'h392;
        15'h117B: data = 12'h4A5;
        15'h117C: data = 12'h5A7;
        15'h117D: data = 12'h6B0;
        15'h117E: data = 12'h7A6;
        15'h117F: data = 12'h0D6;
        15'h1180: data = 12'h1B5;
        15'h1181: data = 12'h28C;
        15'h1182: data = 12'h342;
        15'h1183: data = 12'h3F9;
        15'h1184: data = 12'h499;
        15'h1185: data = 12'h519;
        15'h1186: data = 12'h583;
        15'h1187: data = 12'h5E7;
        15'h1188: data = 12'h626;
        15'h1189: data = 12'h665;
        15'h118A: data = 12'h68C;
        15'h118B: data = 12'h68D;
        15'h118C: data = 12'h693;
        15'h118D: data = 12'h50D;
        15'h118E: data = 12'h63B;
        15'h118F: data = 12'h5E2;
        15'h1190: data = 12'h575;
        15'h1191: data = 12'h504;
        15'h1192: data = 12'h471;
        15'h1193: data = 12'h3D1;
        15'h1194: data = 12'h320;
        15'h1195: data = 12'h266;
        15'h1196: data = 12'h192;
        15'h1197: data = 12'h0B5;
        15'h1198: data = 12'h791;
        15'h1199: data = 12'h69E;
        15'h119A: data = 12'h59A;
        15'h119B: data = 12'h496;
        15'h119C: data = 12'h377;
        15'h119D: data = 12'h25E;
        15'h119E: data = 12'h13C;
        15'h119F: data = 12'h016;
        15'h11A0: data = 12'h6A6;
        15'h11A1: data = 12'h57B;
        15'h11A2: data = 12'h467;
        15'h11A3: data = 12'h348;
        15'h11A4: data = 12'h23D;
        15'h11A5: data = 12'h12C;
        15'h11A6: data = 12'h036;
        15'h11A7: data = 12'h704;
        15'h11A8: data = 12'h615;
        15'h11A9: data = 12'h530;
        15'h11AA: data = 12'h463;
        15'h11AB: data = 12'h393;
        15'h11AC: data = 12'h50D;
        15'h11AD: data = 12'h22F;
        15'h11AE: data = 12'h196;
        15'h11AF: data = 12'h10D;
        15'h11B0: data = 12'h0B6;
        15'h11B1: data = 12'h05F;
        15'h11B2: data = 12'h7C3;
        15'h11B3: data = 12'h782;
        15'h11B4: data = 12'h778;
        15'h11B5: data = 12'h761;
        15'h11B6: data = 12'h781;
        15'h11B7: data = 12'h7A3;
        15'h11B8: data = 12'h7E5;
        15'h11B9: data = 12'h093;
        15'h11BA: data = 12'h0FA;
        15'h11BB: data = 12'h16E;
        15'h11BC: data = 12'h205;
        15'h11BD: data = 12'h2AD;
        15'h11BE: data = 12'h366;
        15'h11BF: data = 12'h437;
        15'h11C0: data = 12'h507;
        15'h11C1: data = 12'h5ED;
        15'h11C2: data = 12'h6D8;
        15'h11C3: data = 12'h7CF;
        15'h11C4: data = 12'h0FA;
        15'h11C5: data = 12'h201;
        15'h11C6: data = 12'h30B;
        15'h11C7: data = 12'h428;
        15'h11C8: data = 12'h53F;
        15'h11C9: data = 12'h66C;
        15'h11CA: data = 12'h798;
        15'h11CB: data = 12'h50D;
        15'h11CC: data = 12'h21F;
        15'h11CD: data = 12'h343;
        15'h11CE: data = 12'h455;
        15'h11CF: data = 12'h55A;
        15'h11D0: data = 12'h659;
        15'h11D1: data = 12'h752;
        15'h11D2: data = 12'h279;
        15'h11D3: data = 12'h168;
        15'h11D4: data = 12'h23D;
        15'h11D5: data = 12'h306;
        15'h11D6: data = 12'h3C4;
        15'h11D7: data = 12'h464;
        15'h11D8: data = 12'h4F4;
        15'h11D9: data = 12'h568;
        15'h11DA: data = 12'h5CC;
        15'h11DB: data = 12'h607;
        15'h11DC: data = 12'h647;
        15'h11DD: data = 12'h678;
        15'h11DE: data = 12'h683;
        15'h11DF: data = 12'h686;
        15'h11E0: data = 12'h66D;
        15'h11E1: data = 12'h641;
        15'h11E2: data = 12'h5F7;
        15'h11E3: data = 12'h59D;
        15'h11E4: data = 12'h53A;
        15'h11E5: data = 12'h4AA;
        15'h11E6: data = 12'h412;
        15'h11E7: data = 12'h35F;
        15'h11E8: data = 12'h2A4;
        15'h11E9: data = 12'h1D5;
        15'h11EA: data = 12'h50D;
        15'h11EB: data = 12'h056;
        15'h11EC: data = 12'h6E3;
        15'h11ED: data = 12'h5ED;
        15'h11EE: data = 12'h4E2;
        15'h11EF: data = 12'h3D3;
        15'h11F0: data = 12'h2B7;
        15'h11F1: data = 12'h19F;
        15'h11F2: data = 12'h082;
        15'h11F3: data = 12'h708;
        15'h11F4: data = 12'h5ED;
        15'h11F5: data = 12'h4CE;
        15'h11F6: data = 12'h3A3;
        15'h11F7: data = 12'h291;
        15'h11F8: data = 12'h17A;
        15'h11F9: data = 12'h07F;
        15'h11FA: data = 12'h74B;
        15'h11FB: data = 12'h665;
        15'h11FC: data = 12'h577;
        15'h11FD: data = 12'h4A5;
        15'h11FE: data = 12'h3D7;
        15'h11FF: data = 12'h31C;
        15'h1200: data = 12'h26C;
        15'h1201: data = 12'h1D5;
        15'h1202: data = 12'h13D;
        15'h1203: data = 12'h0D8;
        15'h1204: data = 12'h076;
        15'h1205: data = 12'h025;
        15'h1206: data = 12'h797;
        15'h1207: data = 12'h77A;
        15'h1208: data = 12'h75D;
        15'h1209: data = 12'h50D;
        15'h120A: data = 12'h7A5;
        15'h120B: data = 12'h7E5;
        15'h120C: data = 12'h741;
        15'h120D: data = 12'h0E0;
        15'h120E: data = 12'h14D;
        15'h120F: data = 12'h1D0;
        15'h1210: data = 12'h26B;
        15'h1211: data = 12'h321;
        15'h1212: data = 12'h3E3;
        15'h1213: data = 12'h4BA;
        15'h1214: data = 12'h598;
        15'h1215: data = 12'h689;
        15'h1216: data = 12'h77D;
        15'h1217: data = 12'h0AE;
        15'h1218: data = 12'h1AC;
        15'h1219: data = 12'h2C3;
        15'h121A: data = 12'h3CF;
        15'h121B: data = 12'h4EB;
        15'h121C: data = 12'h607;
        15'h121D: data = 12'h720;
        15'h121E: data = 12'h3BA;
        15'h121F: data = 12'h1BC;
        15'h1220: data = 12'h2E2;
        15'h1221: data = 12'h401;
        15'h1222: data = 12'h510;
        15'h1223: data = 12'h616;
        15'h1224: data = 12'h70E;
        15'h1225: data = 12'h7F8;
        15'h1226: data = 12'h116;
        15'h1227: data = 12'h1E8;
        15'h1228: data = 12'h50D;
        15'h1229: data = 12'h373;
        15'h122A: data = 12'h423;
        15'h122B: data = 12'h4BD;
        15'h122C: data = 12'h547;
        15'h122D: data = 12'h5AD;
        15'h122E: data = 12'h5FC;
        15'h122F: data = 12'h64A;
        15'h1230: data = 12'h669;
        15'h1231: data = 12'h683;
        15'h1232: data = 12'h682;
        15'h1233: data = 12'h664;
        15'h1234: data = 12'h646;
        15'h1235: data = 12'h606;
        15'h1236: data = 12'h5BC;
        15'h1237: data = 12'h559;
        15'h1238: data = 12'h4DD;
        15'h1239: data = 12'h44C;
        15'h123A: data = 12'h3A1;
        15'h123B: data = 12'h2ED;
        15'h123C: data = 12'h21B;
        15'h123D: data = 12'h148;
        15'h123E: data = 12'h063;
        15'h123F: data = 12'h72F;
        15'h1240: data = 12'h633;
        15'h1241: data = 12'h534;
        15'h1242: data = 12'h424;
        15'h1243: data = 12'h31B;
        15'h1244: data = 12'h1FE;
        15'h1245: data = 12'h0DC;
        15'h1246: data = 12'h771;
        15'h1247: data = 12'h50D;
        15'h1248: data = 12'h52F;
        15'h1249: data = 12'h414;
        15'h124A: data = 12'h2F1;
        15'h124B: data = 12'h1D8;
        15'h124C: data = 12'h0CE;
        15'h124D: data = 12'h7A1;
        15'h124E: data = 12'h6A6;
        15'h124F: data = 12'h5C1;
        15'h1250: data = 12'h4EB;
        15'h1251: data = 12'h419;
        15'h1252: data = 12'h358;
        15'h1253: data = 12'h2A0;
        15'h1254: data = 12'h1FE;
        15'h1255: data = 12'h175;
        15'h1256: data = 12'h100;
        15'h1257: data = 12'h09A;
        15'h1258: data = 12'h039;
        15'h1259: data = 12'h793;
        15'h125A: data = 12'h772;
        15'h125B: data = 12'h755;
        15'h125C: data = 12'h778;
        15'h125D: data = 12'h77E;
        15'h125E: data = 12'h7C0;
        15'h125F: data = 12'h809;
        15'h1260: data = 12'h0C4;
        15'h1261: data = 12'h12C;
        15'h1262: data = 12'h1B1;
        15'h1263: data = 12'h245;
        15'h1264: data = 12'h2E8;
        15'h1265: data = 12'h39B;
        15'h1266: data = 12'h50D;
        15'h1267: data = 12'h541;
        15'h1268: data = 12'h632;
        15'h1269: data = 12'h724;
        15'h126A: data = 12'h828;
        15'h126B: data = 12'h15D;
        15'h126C: data = 12'h26A;
        15'h126D: data = 12'h380;
        15'h126E: data = 12'h495;
        15'h126F: data = 12'h5A6;
        15'h1270: data = 12'h6D0;
        15'h1271: data = 12'h7E8;
        15'h1272: data = 12'h153;
        15'h1273: data = 12'h279;
        15'h1274: data = 12'h394;
        15'h1275: data = 12'h4B3;
        15'h1276: data = 12'h5B7;
        15'h1277: data = 12'h6C4;
        15'h1278: data = 12'h7B1;
        15'h1279: data = 12'h0D9;
        15'h127A: data = 12'h1B2;
        15'h127B: data = 12'h27F;
        15'h127C: data = 12'h332;
        15'h127D: data = 12'h3ED;
        15'h127E: data = 12'h48B;
        15'h127F: data = 12'h514;
        15'h1280: data = 12'h588;
        15'h1281: data = 12'h5F6;
        15'h1282: data = 12'h639;
        15'h1283: data = 12'h679;
        15'h1284: data = 12'h694;
        15'h1285: data = 12'h50D;
        15'h1286: data = 12'h68A;
        15'h1287: data = 12'h660;
        15'h1288: data = 12'h626;
        15'h1289: data = 12'h5D5;
        15'h128A: data = 12'h56D;
        15'h128B: data = 12'h508;
        15'h128C: data = 12'h47C;
        15'h128D: data = 12'h3E2;
        15'h128E: data = 12'h333;
        15'h128F: data = 12'h26F;
        15'h1290: data = 12'h19A;
        15'h1291: data = 12'h0BD;
        15'h1292: data = 12'h78D;
        15'h1293: data = 12'h691;
        15'h1294: data = 12'h589;
        15'h1295: data = 12'h47B;
        15'h1296: data = 12'h364;
        15'h1297: data = 12'h24E;
        15'h1298: data = 12'h139;
        15'h1299: data = 12'h1E9;
        15'h129A: data = 12'h6B8;
        15'h129B: data = 12'h590;
        15'h129C: data = 12'h478;
        15'h129D: data = 12'h357;
        15'h129E: data = 12'h23E;
        15'h129F: data = 12'h120;
        15'h12A0: data = 12'h01E;
        15'h12A1: data = 12'h6F1;
        15'h12A2: data = 12'h603;
        15'h12A3: data = 12'h524;
        15'h12A4: data = 12'h50D;
        15'h12A5: data = 12'h392;
        15'h12A6: data = 12'h2E1;
        15'h12A7: data = 12'h236;
        15'h12A8: data = 12'h1A3;
        15'h12A9: data = 12'h11C;
        15'h12AA: data = 12'h0BF;
        15'h12AB: data = 12'h061;
        15'h12AC: data = 12'h7A7;
        15'h12AD: data = 12'h771;
        15'h12AE: data = 12'h765;
        15'h12AF: data = 12'h751;
        15'h12B0: data = 12'h774;
        15'h12B1: data = 12'h79E;
        15'h12B2: data = 12'h7E7;
        15'h12B3: data = 12'h0C8;
        15'h12B4: data = 12'h10B;
        15'h12B5: data = 12'h180;
        15'h12B6: data = 12'h212;
        15'h12B7: data = 12'h2B5;
        15'h12B8: data = 12'h363;
        15'h12B9: data = 12'h423;
        15'h12BA: data = 12'h4F6;
        15'h12BB: data = 12'h5D9;
        15'h12BC: data = 12'h6CE;
        15'h12BD: data = 12'h7CC;
        15'h12BE: data = 12'h105;
        15'h12BF: data = 12'h20C;
        15'h12C0: data = 12'h31B;
        15'h12C1: data = 12'h43E;
        15'h12C2: data = 12'h54F;
        15'h12C3: data = 12'h50D;
        15'h12C4: data = 12'h78C;
        15'h12C5: data = 12'h0F4;
        15'h12C6: data = 12'h20D;
        15'h12C7: data = 12'h332;
        15'h12C8: data = 12'h44B;
        15'h12C9: data = 12'h55D;
        15'h12CA: data = 12'h669;
        15'h12CB: data = 12'h763;
        15'h12CC: data = 12'h57B;
        15'h12CD: data = 12'h171;
        15'h12CE: data = 12'h23F;
        15'h12CF: data = 12'h2FC;
        15'h12D0: data = 12'h3AD;
        15'h12D1: data = 12'h452;
        15'h12D2: data = 12'h4E3;
        15'h12D3: data = 12'h55A;
        15'h12D4: data = 12'h5CF;
        15'h12D5: data = 12'h611;
        15'h12D6: data = 12'h657;
        15'h12D7: data = 12'h685;
        15'h12D8: data = 12'h691;
        15'h12D9: data = 12'h693;
        15'h12DA: data = 12'h66A;
        15'h12DB: data = 12'h62D;
        15'h12DC: data = 12'h5E2;
        15'h12DD: data = 12'h58B;
        15'h12DE: data = 12'h528;
        15'h12DF: data = 12'h49E;
        15'h12E0: data = 12'h414;
        15'h12E1: data = 12'h369;
        15'h12E2: data = 12'h50D;
        15'h12E3: data = 12'h1E5;
        15'h12E4: data = 12'h109;
        15'h12E5: data = 12'h01F;
        15'h12E6: data = 12'h6E6;
        15'h12E7: data = 12'h5E7;
        15'h12E8: data = 12'h4D2;
        15'h12E9: data = 12'h3C1;
        15'h12EA: data = 12'h2AA;
        15'h12EB: data = 12'h18E;
        15'h12EC: data = 12'h07A;
        15'h12ED: data = 12'h704;
        15'h12EE: data = 12'h5F5;
        15'h12EF: data = 12'h4DD;
        15'h12F0: data = 12'h3B6;
        15'h12F1: data = 12'h2A0;
        15'h12F2: data = 12'h187;
        15'h12F3: data = 12'h086;
        15'h12F4: data = 12'h744;
        15'h12F5: data = 12'h65D;
        15'h12F6: data = 12'h569;
        15'h12F7: data = 12'h49A;
        15'h12F8: data = 12'h3CA;
        15'h12F9: data = 12'h30A;
        15'h12FA: data = 12'h26B;
        15'h12FB: data = 12'h1D5;
        15'h12FC: data = 12'h145;
        15'h12FD: data = 12'h0E6;
        15'h12FE: data = 12'h08A;
        15'h12FF: data = 12'h034;
        15'h1300: data = 12'h79A;
        15'h1301: data = 12'h50D;
        15'h1302: data = 12'h753;
        15'h1303: data = 12'h773;
        15'h1304: data = 12'h793;
        15'h1305: data = 12'h7D4;
        15'h1306: data = 12'h31F;
        15'h1307: data = 12'h0E1;
        15'h1308: data = 12'h159;
        15'h1309: data = 12'h1E2;
        15'h130A: data = 12'h27F;
        15'h130B: data = 12'h333;
        15'h130C: data = 12'h3EC;
        15'h130D: data = 12'h4B6;
        15'h130E: data = 12'h58B;
        15'h130F: data = 12'h676;
        15'h1310: data = 12'h76C;
        15'h1311: data = 12'h0FF;
        15'h1312: data = 12'h1A7;
        15'h1313: data = 12'h2CD;
        15'h1314: data = 12'h3DF;
        15'h1315: data = 12'h502;
        15'h1316: data = 12'h611;
        15'h1317: data = 12'h725;
        15'h1318: data = 12'h4E2;
        15'h1319: data = 12'h1B2;
        15'h131A: data = 12'h2CE;
        15'h131B: data = 12'h3EC;
        15'h131C: data = 12'h504;
        15'h131D: data = 12'h612;
        15'h131E: data = 12'h711;
        15'h131F: data = 12'h801;
        15'h1320: data = 12'h50D;
        15'h1321: data = 12'h1FB;
        15'h1322: data = 12'h2C6;
        15'h1323: data = 12'h37B;
        15'h1324: data = 12'h41A;
        15'h1325: data = 12'h4AD;
        15'h1326: data = 12'h535;
        15'h1327: data = 12'h5A3;
        15'h1328: data = 12'h5F2;
        15'h1329: data = 12'h64E;
        15'h132A: data = 12'h678;
        15'h132B: data = 12'h697;
        15'h132C: data = 12'h695;
        15'h132D: data = 12'h673;
        15'h132E: data = 12'h64B;
        15'h132F: data = 12'h601;
        15'h1330: data = 12'h5AD;
        15'h1331: data = 12'h543;
        15'h1332: data = 12'h4CC;
        15'h1333: data = 12'h445;
        15'h1334: data = 12'h39F;
        15'h1335: data = 12'h2F0;
        15'h1336: data = 12'h22B;
        15'h1337: data = 12'h14F;
        15'h1338: data = 12'h06A;
        15'h1339: data = 12'h740;
        15'h133A: data = 12'h63D;
        15'h133B: data = 12'h535;
        15'h133C: data = 12'h41C;
        15'h133D: data = 12'h30D;
        15'h133E: data = 12'h1EA;
        15'h133F: data = 12'h50D;
        15'h1340: data = 12'h76B;
        15'h1341: data = 12'h648;
        15'h1342: data = 12'h52D;
        15'h1343: data = 12'h41B;
        15'h1344: data = 12'h2FE;
        15'h1345: data = 12'h1E9;
        15'h1346: data = 12'h0DC;
        15'h1347: data = 12'h78B;
        15'h1348: data = 12'h6AA;
        15'h1349: data = 12'h5B7;
        15'h134A: data = 12'h4E0;
        15'h134B: data = 12'h40B;
        15'h134C: data = 12'h348;
        15'h134D: data = 12'h29C;
        15'h134E: data = 12'h1FD;
        15'h134F: data = 12'h175;
        15'h1350: data = 12'h103;
        15'h1351: data = 12'h0A0;
        15'h1352: data = 12'h048;
        15'h1353: data = 12'h7A0;
        15'h1354: data = 12'h77F;
        15'h1355: data = 12'h75B;
        15'h1356: data = 12'h774;
        15'h1357: data = 12'h778;
        15'h1358: data = 12'h7B2;
        15'h1359: data = 12'h7F7;
        15'h135A: data = 12'h0BC;
        15'h135B: data = 12'h125;
        15'h135C: data = 12'h1B5;
        15'h135D: data = 12'h250;
        15'h135E: data = 12'h50D;
        15'h135F: data = 12'h3AD;
        15'h1360: data = 12'h47B;
        15'h1361: data = 12'h53D;
        15'h1362: data = 12'h62A;
        15'h1363: data = 12'h717;
        15'h1364: data = 12'h81C;
        15'h1365: data = 12'h154;
        15'h1366: data = 12'h269;
        15'h1367: data = 12'h385;
        15'h1368: data = 12'h4A1;
        15'h1369: data = 12'h5B3;
        15'h136A: data = 12'h6DE;
        15'h136B: data = 12'h7F2;
        15'h136C: data = 12'h155;
        15'h136D: data = 12'h276;
        15'h136E: data = 12'h38C;
        15'h136F: data = 12'h4A7;
        15'h1370: data = 12'h5B1;
        15'h1371: data = 12'h6BE;
        15'h1372: data = 12'h7B6;
        15'h1373: data = 12'h0E0;
        15'h1374: data = 12'h1BF;
        15'h1375: data = 12'h28C;
        15'h1376: data = 12'h340;
        15'h1377: data = 12'h3F1;
        15'h1378: data = 12'h48B;
        15'h1379: data = 12'h510;
        15'h137A: data = 12'h580;
        15'h137B: data = 12'h5EE;
        15'h137C: data = 12'h637;
        15'h137D: data = 12'h50D;
        15'h137E: data = 12'h69B;
        15'h137F: data = 12'h69B;
        15'h1380: data = 12'h698;
        15'h1381: data = 12'h66F;
        15'h1382: data = 12'h632;
        15'h1383: data = 12'h5D5;
        15'h1384: data = 12'h568;
        15'h1385: data = 12'h4FE;
        15'h1386: data = 12'h470;
        15'h1387: data = 12'h3DB;
        15'h1388: data = 12'h32F;
        15'h1389: data = 12'h270;
        15'h138A: data = 12'h1A4;
        15'h138B: data = 12'h0C3;
        15'h138C: data = 12'h78C;
        15'h138D: data = 12'h699;
        15'h138E: data = 12'h58F;
        15'h138F: data = 12'h483;
        15'h1390: data = 12'h365;
        15'h1391: data = 12'h24C;
        15'h1392: data = 12'h133;
        15'h1393: data = 12'h062;
        15'h1394: data = 12'h6AD;
        15'h1395: data = 12'h589;
        15'h1396: data = 12'h476;
        15'h1397: data = 12'h35A;
        15'h1398: data = 12'h245;
        15'h1399: data = 12'h12F;
        15'h139A: data = 12'h031;
        15'h139B: data = 12'h701;
        15'h139C: data = 12'h50D;
        15'h139D: data = 12'h524;
        15'h139E: data = 12'h455;
        15'h139F: data = 12'h388;
        15'h13A0: data = 12'h2D4;
        15'h13A1: data = 12'h22F;
        15'h13A2: data = 12'h19E;
        15'h13A3: data = 12'h11D;
        15'h13A4: data = 12'h0C8;
        15'h13A5: data = 12'h068;
        15'h13A6: data = 12'h758;
        15'h13A7: data = 12'h77F;
        15'h13A8: data = 12'h76F;
        15'h13A9: data = 12'h757;
        15'h13AA: data = 12'h772;
        15'h13AB: data = 12'h798;
        15'h13AC: data = 12'h7E2;
        15'h13AD: data = 12'h099;
        15'h13AE: data = 12'h104;
        15'h13AF: data = 12'h17E;
        15'h13B0: data = 12'h216;
        15'h13B1: data = 12'h2BB;
        15'h13B2: data = 12'h372;
        15'h13B3: data = 12'h435;
        15'h13B4: data = 12'h501;
        15'h13B5: data = 12'h5DC;
        15'h13B6: data = 12'h6CD;
        15'h13B7: data = 12'h7C2;
        15'h13B8: data = 12'h0F8;
        15'h13B9: data = 12'h209;
        15'h13BA: data = 12'h31A;
        15'h13BB: data = 12'h50D;
        15'h13BC: data = 12'h556;
        15'h13BD: data = 12'h67D;
        15'h13BE: data = 12'h79A;
        15'h13BF: data = 12'h0FD;
        15'h13C0: data = 12'h210;
        15'h13C1: data = 12'h330;
        15'h13C2: data = 12'h446;
        15'h13C3: data = 12'h559;
        15'h13C4: data = 12'h660;
        15'h13C5: data = 12'h765;
        15'h13C6: data = 12'h48C;
        15'h13C7: data = 12'h176;
        15'h13C8: data = 12'h246;
        15'h13C9: data = 12'h302;
        15'h13CA: data = 12'h3B2;
        15'h13CB: data = 12'h44F;
        15'h13CC: data = 12'h4E3;
        15'h13CD: data = 12'h558;
        15'h13CE: data = 12'h5C9;
        15'h13CF: data = 12'h613;
        15'h13D0: data = 12'h652;
        15'h13D1: data = 12'h68C;
        15'h13D2: data = 12'h699;
        15'h13D3: data = 12'h69A;
        15'h13D4: data = 12'h675;
        15'h13D5: data = 12'h634;
        15'h13D6: data = 12'h5E4;
        15'h13D7: data = 12'h58A;
        15'h13D8: data = 12'h52B;
        15'h13D9: data = 12'h49B;
        15'h13DA: data = 12'h50D;
        15'h13DB: data = 12'h364;
        15'h13DC: data = 12'h2AE;
        15'h13DD: data = 12'h1E6;
        15'h13DE: data = 12'h110;
        15'h13DF: data = 12'h023;
        15'h13E0: data = 12'h6F1;
        15'h13E1: data = 12'h5EF;
        15'h13E2: data = 12'h4DD;
        15'h13E3: data = 12'h3C5;
        15'h13E4: data = 12'h2A8;
        15'h13E5: data = 12'h18D;
        15'h13E6: data = 12'h070;
        15'h13E7: data = 12'h6FC;
        15'h13E8: data = 12'h5EA;
        15'h13E9: data = 12'h4D9;
        15'h13EA: data = 12'h3B7;
        15'h13EB: data = 12'h2A7;
        15'h13EC: data = 12'h18F;
        15'h13ED: data = 12'h08B;
        15'h13EE: data = 12'h74A;
        15'h13EF: data = 12'h65C;
        15'h13F0: data = 12'h569;
        15'h13F1: data = 12'h491;
        15'h13F2: data = 12'h3C6;
        15'h13F3: data = 12'h30D;
        15'h13F4: data = 12'h267;
        15'h13F5: data = 12'h1D1;
        15'h13F6: data = 12'h141;
        15'h13F7: data = 12'h0E5;
        15'h13F8: data = 12'h088;
        15'h13F9: data = 12'h50D;
        15'h13FA: data = 12'h7A4;
        15'h13FB: data = 12'h77E;
        15'h13FC: data = 12'h75B;
        15'h13FD: data = 12'h776;
        15'h13FE: data = 12'h795;
        15'h13FF: data = 12'h7D3;
        15'h1400: data = 12'h289;
        15'h1401: data = 12'h0E2;
        15'h1402: data = 12'h155;
        15'h1403: data = 12'h1E2;
        15'h1404: data = 12'h27F;
        15'h1405: data = 12'h339;
        15'h1406: data = 12'h3F5;
        15'h1407: data = 12'h4C1;
        15'h1408: data = 12'h590;
        15'h1409: data = 12'h67C;
        15'h140A: data = 12'h76B;
        15'h140B: data = 12'h107;
        15'h140C: data = 12'h1A5;
        15'h140D: data = 12'h2C8;
        15'h140E: data = 12'h3DD;
        15'h140F: data = 12'h502;
        15'h1410: data = 12'h61E;
        15'h1411: data = 12'h731;
        15'h1412: data = 12'h55A;
        15'h1413: data = 12'h1B7;
        15'h1414: data = 12'h2D3;
        15'h1415: data = 12'h3EF;
        15'h1416: data = 12'h500;
        15'h1417: data = 12'h60B;
        15'h1418: data = 12'h50D;
        15'h1419: data = 12'h804;
        15'h141A: data = 12'h12A;
        15'h141B: data = 12'h1FC;
        15'h141C: data = 12'h2C9;
        15'h141D: data = 12'h37E;
        15'h141E: data = 12'h422;
        15'h141F: data = 12'h4AE;
        15'h1420: data = 12'h532;
        15'h1421: data = 12'h5A4;
        15'h1422: data = 12'h5F1;
        15'h1423: data = 12'h64E;
        15'h1424: data = 12'h670;
        15'h1425: data = 12'h69A;
        15'h1426: data = 12'h695;
        15'h1427: data = 12'h676;
        15'h1428: data = 12'h653;
        15'h1429: data = 12'h612;
        15'h142A: data = 12'h5B6;
        15'h142B: data = 12'h54D;
        15'h142C: data = 12'h4C7;
        15'h142D: data = 12'h43E;
        15'h142E: data = 12'h392;
        15'h142F: data = 12'h2E6;
        15'h1430: data = 12'h220;
        15'h1431: data = 12'h14D;
        15'h1432: data = 12'h073;
        15'h1433: data = 12'h743;
        15'h1434: data = 12'h641;
        15'h1435: data = 12'h53D;
        15'h1436: data = 12'h429;
        15'h1437: data = 12'h50D;
        15'h1438: data = 12'h1EF;
        15'h1439: data = 12'h0D2;
        15'h143A: data = 12'h768;
        15'h143B: data = 12'h63F;
        15'h143C: data = 12'h524;
        15'h143D: data = 12'h414;
        15'h143E: data = 12'h2FE;
        15'h143F: data = 12'h1E9;
        15'h1440: data = 12'h0DE;
        15'h1441: data = 12'h789;
        15'h1442: data = 12'h6AF;
        15'h1443: data = 12'h5C1;
        15'h1444: data = 12'h4E5;
        15'h1445: data = 12'h409;
        15'h1446: data = 12'h347;
        15'h1447: data = 12'h293;
        15'h1448: data = 12'h1F2;
        15'h1449: data = 12'h171;
        15'h144A: data = 12'h103;
        15'h144B: data = 12'h0A2;
        15'h144C: data = 12'h047;
        15'h144D: data = 12'h7A3;
        15'h144E: data = 12'h784;
        15'h144F: data = 12'h75D;
        15'h1450: data = 12'h77C;
        15'h1451: data = 12'h779;
        15'h1452: data = 12'h7B1;
        15'h1453: data = 12'h7F4;
        15'h1454: data = 12'h0B5;
        15'h1455: data = 12'h11F;
        15'h1456: data = 12'h50D;
        15'h1457: data = 12'h24C;
        15'h1458: data = 12'h2F7;
        15'h1459: data = 12'h3B2;
        15'h145A: data = 12'h481;
        15'h145B: data = 12'h54A;
        15'h145C: data = 12'h631;
        15'h145D: data = 12'h714;
        15'h145E: data = 12'h818;
        15'h145F: data = 12'h14D;
        15'h1460: data = 12'h25D;
        15'h1461: data = 12'h37F;
        15'h1462: data = 12'h49D;
        15'h1463: data = 12'h5B7;
        15'h1464: data = 12'h6E3;
        15'h1465: data = 12'h7F8;
        15'h1466: data = 12'h15E;
        15'h1467: data = 12'h279;
        15'h1468: data = 12'h38B;
        15'h1469: data = 12'h4A1;
        15'h146A: data = 12'h5A8;
        15'h146B: data = 12'h6BC;
        15'h146C: data = 12'h7AF;
        15'h146D: data = 12'h0E4;
        15'h146E: data = 12'h1C1;
        15'h146F: data = 12'h292;
        15'h1470: data = 12'h344;
        15'h1471: data = 12'h3F4;
        15'h1472: data = 12'h48B;
        15'h1473: data = 12'h50C;
        15'h1474: data = 12'h578;
        15'h1475: data = 12'h50D;
        15'h1476: data = 12'h630;
        15'h1477: data = 12'h672;
        15'h1478: data = 12'h693;
        15'h1479: data = 12'h697;
        15'h147A: data = 12'h694;
        15'h147B: data = 12'h66D;
        15'h147C: data = 12'h636;
        15'h147D: data = 12'h5D2;
        15'h147E: data = 12'h567;
        15'h147F: data = 12'h4F8;
        15'h1480: data = 12'h46E;
        15'h1481: data = 12'h3CF;
        15'h1482: data = 12'h328;
        15'h1483: data = 12'h268;
        15'h1484: data = 12'h19A;
        15'h1485: data = 12'h0C3;
        15'h1486: data = 12'h792;
        15'h1487: data = 12'h69B;
        15'h1488: data = 12'h594;
        15'h1489: data = 12'h489;
        15'h148A: data = 12'h365;
        15'h148B: data = 12'h24B;
        15'h148C: data = 12'h12E;
        15'h148D: data = 12'h061;
        15'h148E: data = 12'h6A4;
        15'h148F: data = 12'h587;
        15'h1490: data = 12'h473;
        15'h1491: data = 12'h359;
        15'h1492: data = 12'h245;
        15'h1493: data = 12'h132;
        15'h1494: data = 12'h50D;
        15'h1495: data = 12'h703;
        15'h1496: data = 12'h60C;
        15'h1497: data = 12'h523;
        15'h1498: data = 12'h453;
        15'h1499: data = 12'h387;
        15'h149A: data = 12'h2CD;
        15'h149B: data = 12'h22A;
        15'h149C: data = 12'h199;
        15'h149D: data = 12'h117;
        15'h149E: data = 12'h0BF;
        15'h149F: data = 12'h066;
        15'h14A0: data = 12'h777;
        15'h14A1: data = 12'h784;
        15'h14A2: data = 12'h773;
        15'h14A3: data = 12'h75B;
        15'h14A4: data = 12'h775;
        15'h14A5: data = 12'h799;
        15'h14A6: data = 12'h7DE;
        15'h14A7: data = 12'h095;
        15'h14A8: data = 12'h101;
        15'h14A9: data = 12'h17C;
        15'h14AA: data = 12'h216;
        15'h14AB: data = 12'h2BB;
        15'h14AC: data = 12'h374;
        15'h14AD: data = 12'h438;
        15'h14AE: data = 12'h502;
        15'h14AF: data = 12'h5E2;
        15'h14B0: data = 12'h6D0;
        15'h14B1: data = 12'h7C5;
        15'h14B2: data = 12'h0F7;
        15'h14B3: data = 12'h50D;
        15'h14B4: data = 12'h318;
        15'h14B5: data = 12'h441;
        15'h14B6: data = 12'h557;
        15'h14B7: data = 12'h678;
        15'h14B8: data = 12'h79A;
        15'h14B9: data = 12'h100;
        15'h14BA: data = 12'h216;
        15'h14BB: data = 12'h333;
        15'h14BC: data = 12'h444;
        15'h14BD: data = 12'h557;
        15'h14BE: data = 12'h65F;
        15'h14BF: data = 12'h761;
        15'h14C0: data = 12'h1D7;
        15'h14C1: data = 12'h176;
        15'h14C2: data = 12'h247;
        15'h14C3: data = 12'h309;
        15'h14C4: data = 12'h3B9;
        15'h14C5: data = 12'h452;
        15'h14C6: data = 12'h4E0;
        15'h14C7: data = 12'h55A;
        15'h14C8: data = 12'h5C6;
        15'h14C9: data = 12'h60A;
        15'h14CA: data = 12'h64F;
        15'h14CB: data = 12'h68B;
        15'h14CC: data = 12'h694;
        15'h14CD: data = 12'h693;
        15'h14CE: data = 12'h677;
        15'h14CF: data = 12'h639;
        15'h14D0: data = 12'h5E9;
        15'h14D1: data = 12'h58C;
        15'h14D2: data = 12'h50D;
        15'h14D3: data = 12'h49A;
        15'h14D4: data = 12'h409;
        15'h14D5: data = 12'h35B;
        15'h14D6: data = 12'h2A9;
        15'h14D7: data = 12'h1E0;
        15'h14D8: data = 12'h10A;
        15'h14D9: data = 12'h1DF;
        15'h14DA: data = 12'h6F1;
        15'h14DB: data = 12'h5F2;
        15'h14DC: data = 12'h4E0;
        15'h14DD: data = 12'h3C9;
        15'h14DE: data = 12'h2A7;
        15'h14DF: data = 12'h18E;
        15'h14E0: data = 12'h070;
        15'h14E1: data = 12'h6F8;
        15'h14E2: data = 12'h5E4;
        15'h14E3: data = 12'h4D3;
        15'h14E4: data = 12'h3B5;
        15'h14E5: data = 12'h2A5;
        15'h14E6: data = 12'h18F;
        15'h14E7: data = 12'h08B;
        15'h14E8: data = 12'h74B;
        15'h14E9: data = 12'h65D;
        15'h14EA: data = 12'h569;
        15'h14EB: data = 12'h493;
        15'h14EC: data = 12'h3C6;
        15'h14ED: data = 12'h30B;
        15'h14EE: data = 12'h264;
        15'h14EF: data = 12'h1D1;
        15'h14F0: data = 12'h141;
        15'h14F1: data = 12'h50D;
        15'h14F2: data = 12'h084;
        15'h14F3: data = 12'h035;
        15'h14F4: data = 12'h7A5;
        15'h14F5: data = 12'h781;
        15'h14F6: data = 12'h761;
        15'h14F7: data = 12'h77B;
        15'h14F8: data = 12'h793;
        15'h14F9: data = 12'h7D0;
        15'h14FA: data = 12'h370;
        15'h14FB: data = 12'h0D7;
        15'h14FC: data = 12'h14B;
        15'h14FD: data = 12'h1DC;
        15'h14FE: data = 12'h27D;
        15'h14FF: data = 12'h338;
        15'h1500: data = 12'h3F3;
        15'h1501: data = 12'h4C2;
        15'h1502: data = 12'h595;
        15'h1503: data = 12'h67F;
        15'h1504: data = 12'h76A;
        15'h1505: data = 12'h11C;
        15'h1506: data = 12'h1A1;
        15'h1507: data = 12'h2C2;
        15'h1508: data = 12'h3D9;
        15'h1509: data = 12'h4FD;
        15'h150A: data = 12'h61B;
        15'h150B: data = 12'h736;
        15'h150C: data = 12'h5C5;
        15'h150D: data = 12'h1BB;
        15'h150E: data = 12'h2D3;
        15'h150F: data = 12'h3EA;
        15'h1510: data = 12'h50D;
        15'h1511: data = 12'h604;
        15'h1512: data = 12'h707;
        15'h1513: data = 12'h7FF;
        15'h1514: data = 12'h125;
        15'h1515: data = 12'h1F7;
        15'h1516: data = 12'h2CB;
        15'h1517: data = 12'h37F;
        15'h1518: data = 12'h425;
        15'h1519: data = 12'h4B7;
        15'h151A: data = 12'h538;
        15'h151B: data = 12'h59F;
        15'h151C: data = 12'h5ED;
        15'h151D: data = 12'h646;
        15'h151E: data = 12'h66B;
        15'h151F: data = 12'h695;
        15'h1520: data = 12'h699;
        15'h1521: data = 12'h678;
        15'h1522: data = 12'h659;
        15'h1523: data = 12'h616;
        15'h1524: data = 12'h5BA;
        15'h1525: data = 12'h54B;
        15'h1526: data = 12'h4CC;
        15'h1527: data = 12'h43D;
        15'h1528: data = 12'h396;
        15'h1529: data = 12'h2E5;
        15'h152A: data = 12'h222;
        15'h152B: data = 12'h14F;
        15'h152C: data = 12'h070;
        15'h152D: data = 12'h73F;
        15'h152E: data = 12'h642;
        15'h152F: data = 12'h50D;
        15'h1530: data = 12'h429;
        15'h1531: data = 12'h316;
        15'h1532: data = 12'h1F6;
        15'h1533: data = 12'h0D3;
        15'h1534: data = 12'h76A;
        15'h1535: data = 12'h63D;
        15'h1536: data = 12'h521;
        15'h1537: data = 12'h40D;
        15'h1538: data = 12'h2F5;
        15'h1539: data = 12'h1E4;
        15'h153A: data = 12'h0DC;
        15'h153B: data = 12'h75B;
        15'h153C: data = 12'h6B4;
        15'h153D: data = 12'h5C9;
        15'h153E: data = 12'h4E9;
        15'h153F: data = 12'h40C;
        15'h1540: data = 12'h344;
        15'h1541: data = 12'h28E;
        15'h1542: data = 12'h1EE;
        15'h1543: data = 12'h169;
        15'h1544: data = 12'h0F7;
        15'h1545: data = 12'h09B;
        15'h1546: data = 12'h041;
        15'h1547: data = 12'h7A3;
        15'h1548: data = 12'h786;
        15'h1549: data = 12'h767;
        15'h154A: data = 12'h77E;
        15'h154B: data = 12'h77C;
        15'h154C: data = 12'h7B1;
        15'h154D: data = 12'h7EE;
        15'h154E: data = 12'h50D;
        15'h154F: data = 12'h11C;
        15'h1550: data = 12'h1AB;
        15'h1551: data = 12'h248;
        15'h1552: data = 12'h2F1;
        15'h1553: data = 12'h3B0;
        15'h1554: data = 12'h481;
        15'h1555: data = 12'h54C;
        15'h1556: data = 12'h636;
        15'h1557: data = 12'h721;
        15'h1558: data = 12'h819;
        15'h1559: data = 12'h14D;
        15'h155A: data = 12'h25A;
        15'h155B: data = 12'h375;
        15'h155C: data = 12'h494;
        15'h155D: data = 12'h5B1;
        15'h155E: data = 12'h6DD;
        15'h155F: data = 12'h7F6;
        15'h1560: data = 12'h164;
        15'h1561: data = 12'h282;
        15'h1562: data = 12'h394;
        15'h1563: data = 12'h4A6;
        15'h1564: data = 12'h5AD;
        15'h1565: data = 12'h6B1;
        15'h1566: data = 12'h7A7;
        15'h1567: data = 12'h0D4;
        15'h1568: data = 12'h1B7;
        15'h1569: data = 12'h28E;
        15'h156A: data = 12'h348;
        15'h156B: data = 12'h3FC;
        15'h156C: data = 12'h49B;
        15'h156D: data = 12'h50D;
        15'h156E: data = 12'h581;
        15'h156F: data = 12'h5E1;
        15'h1570: data = 12'h624;
        15'h1571: data = 12'h669;
        15'h1572: data = 12'h68E;
        15'h1573: data = 12'h690;
        15'h1574: data = 12'h695;
        15'h1575: data = 12'h66F;
        15'h1576: data = 12'h635;
        15'h1577: data = 12'h5DF;
        15'h1578: data = 12'h571;
        15'h1579: data = 12'h501;
        15'h157A: data = 12'h471;
        15'h157B: data = 12'h3D2;
        15'h157C: data = 12'h31F;
        15'h157D: data = 12'h25D;
        15'h157E: data = 12'h191;
        15'h157F: data = 12'h0B0;
        15'h1580: data = 12'h78D;
        15'h1581: data = 12'h69F;
        15'h1582: data = 12'h594;
        15'h1583: data = 12'h490;
        15'h1584: data = 12'h373;
        15'h1585: data = 12'h25A;
        15'h1586: data = 12'h138;
        15'h1587: data = 12'h019;
        15'h1588: data = 12'h6A3;
        15'h1589: data = 12'h57A;
        15'h158A: data = 12'h469;
        15'h158B: data = 12'h34A;
        15'h158C: data = 12'h50D;
        15'h158D: data = 12'h127;
        15'h158E: data = 12'h059;
        15'h158F: data = 12'h700;
        15'h1590: data = 12'h610;
        15'h1591: data = 12'h531;
        15'h1592: data = 12'h461;
        15'h1593: data = 12'h396;
        15'h1594: data = 12'h2DB;
        15'h1595: data = 12'h22F;
        15'h1596: data = 12'h197;
        15'h1597: data = 12'h10D;
        15'h1598: data = 12'h0B4;
        15'h1599: data = 12'h057;
        15'h159A: data = 12'h7BF;
        15'h159B: data = 12'h77F;
        15'h159C: data = 12'h778;
        15'h159D: data = 12'h764;
        15'h159E: data = 12'h783;
        15'h159F: data = 12'h7A8;
        15'h15A0: data = 12'h7E5;
        15'h15A1: data = 12'h091;
        15'h15A2: data = 12'h0FB;
        15'h15A3: data = 12'h16E;
        15'h15A4: data = 12'h205;
        15'h15A5: data = 12'h2AD;
        15'h15A6: data = 12'h367;
        15'h15A7: data = 12'h438;
        15'h15A8: data = 12'h50B;
        15'h15A9: data = 12'h5EB;
        15'h15AA: data = 12'h6DC;
        15'h15AB: data = 12'h50D;
        15'h15AC: data = 12'h0FF;
        15'h15AD: data = 12'h206;
        15'h15AE: data = 12'h30E;
        15'h15AF: data = 12'h432;
        15'h15B0: data = 12'h53F;
        15'h15B1: data = 12'h66B;
        15'h15B2: data = 12'h795;
        15'h15B3: data = 12'h106;
        15'h15B4: data = 12'h220;
        15'h15B5: data = 12'h345;
        15'h15B6: data = 12'h45A;
        15'h15B7: data = 12'h55E;
        15'h15B8: data = 12'h65F;
        15'h15B9: data = 12'h753;
        15'h15BA: data = 12'h2E2;
        15'h15BB: data = 12'h167;
        15'h15BC: data = 12'h23D;
        15'h15BD: data = 12'h30B;
        15'h15BE: data = 12'h3C4;
        15'h15BF: data = 12'h464;
        15'h15C0: data = 12'h4F7;
        15'h15C1: data = 12'h564;
        15'h15C2: data = 12'h5D0;
        15'h15C3: data = 12'h607;
        15'h15C4: data = 12'h645;
        15'h15C5: data = 12'h67A;
        15'h15C6: data = 12'h686;
        15'h15C7: data = 12'h68B;
        15'h15C8: data = 12'h66A;
        15'h15C9: data = 12'h63A;
        15'h15CA: data = 12'h50D;
        15'h15CB: data = 12'h59F;
        15'h15CC: data = 12'h538;
        15'h15CD: data = 12'h4A8;
        15'h15CE: data = 12'h412;
        15'h15CF: data = 12'h35E;
        15'h15D0: data = 12'h29D;
        15'h15D1: data = 12'h1D5;
        15'h15D2: data = 12'h0F8;
        15'h15D3: data = 12'h09C;
        15'h15D4: data = 12'h6DD;
        15'h15D5: data = 12'h5E5;
        15'h15D6: data = 12'h4E0;
        15'h15D7: data = 12'h3D5;
        15'h15D8: data = 12'h2B5;
        15'h15D9: data = 12'h19A;
        15'h15DA: data = 12'h07D;
        15'h15DB: data = 12'h704;
        15'h15DC: data = 12'h5E1;
        15'h15DD: data = 12'h4C8;
        15'h15DE: data = 12'h3A0;
        15'h15DF: data = 12'h290;
        15'h15E0: data = 12'h179;
        15'h15E1: data = 12'h07A;
        15'h15E2: data = 12'h745;
        15'h15E3: data = 12'h65F;
        15'h15E4: data = 12'h573;
        15'h15E5: data = 12'h4A1;
        15'h15E6: data = 12'h3D6;
        15'h15E7: data = 12'h319;
        15'h15E8: data = 12'h271;
        15'h15E9: data = 12'h50D;
        15'h15EA: data = 12'h13C;
        15'h15EB: data = 12'h0D6;
        15'h15EC: data = 12'h073;
        15'h15ED: data = 12'h7BE;
        15'h15EE: data = 12'h792;
        15'h15EF: data = 12'h776;
        15'h15F0: data = 12'h75F;
        15'h15F1: data = 12'h782;
        15'h15F2: data = 12'h7A9;
        15'h15F3: data = 12'h7E2;
        15'h15F4: data = 12'h7A9;
        15'h15F5: data = 12'h0E1;
        15'h15F6: data = 12'h14A;
        15'h15F7: data = 12'h1D1;
        15'h15F8: data = 12'h26E;
        15'h15F9: data = 12'h324;
        15'h15FA: data = 12'h3E4;
        15'h15FB: data = 12'h4B6;
        15'h15FC: data = 12'h598;
        15'h15FD: data = 12'h688;
        15'h15FE: data = 12'h77A;
        15'h15FF: data = 12'h0CE;
        15'h1600: data = 12'h1AE;
        15'h1601: data = 12'h2C3;
        15'h1602: data = 12'h3D4;
        15'h1603: data = 12'h4F2;
        15'h1604: data = 12'h60C;
        15'h1605: data = 12'h726;
        15'h1606: data = 12'h289;
        15'h1607: data = 12'h1C0;
        15'h1608: data = 12'h50D;
        15'h1609: data = 12'h3FE;
        15'h160A: data = 12'h50E;
        15'h160B: data = 12'h618;
        15'h160C: data = 12'h711;
        15'h160D: data = 12'h7FD;
        15'h160E: data = 12'h11A;
        15'h160F: data = 12'h1EB;
        15'h1610: data = 12'h2B7;
        15'h1611: data = 12'h377;
        15'h1612: data = 12'h425;
        15'h1613: data = 12'h4BA;
        15'h1614: data = 12'h54D;
        15'h1615: data = 12'h5B4;
        15'h1616: data = 12'h603;
        15'h1617: data = 12'h654;
        15'h1618: data = 12'h670;
        15'h1619: data = 12'h68B;
        15'h161A: data = 12'h687;
        15'h161B: data = 12'h661;
        15'h161C: data = 12'h641;
        15'h161D: data = 12'h609;
        15'h161E: data = 12'h5BB;
        15'h161F: data = 12'h55A;
        15'h1620: data = 12'h4DC;
        15'h1621: data = 12'h44D;
        15'h1622: data = 12'h3A0;
        15'h1623: data = 12'h2EA;
        15'h1624: data = 12'h21B;
        15'h1625: data = 12'h144;
        15'h1626: data = 12'h062;
        15'h1627: data = 12'h50D;
        15'h1628: data = 12'h62D;
        15'h1629: data = 12'h534;
        15'h162A: data = 12'h420;
        15'h162B: data = 12'h319;
        15'h162C: data = 12'h1FB;
        15'h162D: data = 12'h0E0;
        15'h162E: data = 12'h776;
        15'h162F: data = 12'h64D;
        15'h1630: data = 12'h52B;
        15'h1631: data = 12'h412;
        15'h1632: data = 12'h2F3;
        15'h1633: data = 12'h1D7;
        15'h1634: data = 12'h0CE;
        15'h1635: data = 12'h7A5;
        15'h1636: data = 12'h6A7;
        15'h1637: data = 12'h5BA;
        15'h1638: data = 12'h4E9;
        15'h1639: data = 12'h416;
        15'h163A: data = 12'h354;
        15'h163B: data = 12'h2A2;
        15'h163C: data = 12'h202;
        15'h163D: data = 12'h179;
        15'h163E: data = 12'h102;
        15'h163F: data = 12'h099;
        15'h1640: data = 12'h03B;
        15'h1641: data = 12'h793;
        15'h1642: data = 12'h770;
        15'h1643: data = 12'h753;
        15'h1644: data = 12'h778;
        15'h1645: data = 12'h784;
        15'h1646: data = 12'h50D;
        15'h1647: data = 12'h80A;
        15'h1648: data = 12'h0C5;
        15'h1649: data = 12'h12C;
        15'h164A: data = 12'h1B0;
        15'h164B: data = 12'h249;
        15'h164C: data = 12'h2EA;
        15'h164D: data = 12'h3A2;
        15'h164E: data = 12'h474;
        15'h164F: data = 12'h547;
        15'h1650: data = 12'h633;
        15'h1651: data = 12'h728;
        15'h1652: data = 12'h828;
        15'h1653: data = 12'h161;
        15'h1654: data = 12'h26F;
        15'h1655: data = 12'h384;
        15'h1656: data = 12'h498;
        15'h1657: data = 12'h5AD;
        15'h1658: data = 12'h6D5;
        15'h1659: data = 12'h7E9;
        15'h165A: data = 12'h159;
        15'h165B: data = 12'h280;
        15'h165C: data = 12'h39A;
        15'h165D: data = 12'h4B0;
        15'h165E: data = 12'h5BF;
        15'h165F: data = 12'h6C8;
        15'h1660: data = 12'h7B5;
        15'h1661: data = 12'h0E1;
        15'h1662: data = 12'h1B1;
        15'h1663: data = 12'h27C;
        15'h1664: data = 12'h332;
        15'h1665: data = 12'h50D;
        15'h1666: data = 12'h48B;
        15'h1667: data = 12'h514;
        15'h1668: data = 12'h591;
        15'h1669: data = 12'h5F9;
        15'h166A: data = 12'h639;
        15'h166B: data = 12'h676;
        15'h166C: data = 12'h68F;
        15'h166D: data = 12'h68D;
        15'h166E: data = 12'h684;
        15'h166F: data = 12'h65B;
        15'h1670: data = 12'h627;
        15'h1671: data = 12'h5CF;
        15'h1672: data = 12'h56D;
        15'h1673: data = 12'h503;
        15'h1674: data = 12'h47C;
        15'h1675: data = 12'h3E3;
        15'h1676: data = 12'h330;
        15'h1677: data = 12'h26C;
        15'h1678: data = 12'h197;
        15'h1679: data = 12'h0B6;
        15'h167A: data = 12'h78B;
        15'h167B: data = 12'h68A;
        15'h167C: data = 12'h585;
        15'h167D: data = 12'h47C;
        15'h167E: data = 12'h366;
        15'h167F: data = 12'h252;
        15'h1680: data = 12'h13B;
        15'h1681: data = 12'h218;
        15'h1682: data = 12'h6AF;
        15'h1683: data = 12'h58A;
        15'h1684: data = 12'h50D;
        15'h1685: data = 12'h34F;
        15'h1686: data = 12'h23D;
        15'h1687: data = 12'h122;
        15'h1688: data = 12'h020;
        15'h1689: data = 12'h6F0;
        15'h168A: data = 12'h600;
        15'h168B: data = 12'h523;
        15'h168C: data = 12'h458;
        15'h168D: data = 12'h391;
        15'h168E: data = 12'h2DB;
        15'h168F: data = 12'h23A;
        15'h1690: data = 12'h1A3;
        15'h1691: data = 12'h11B;
        15'h1692: data = 12'h0C0;
        15'h1693: data = 12'h05E;
        15'h1694: data = 12'h7AD;
        15'h1695: data = 12'h774;
        15'h1696: data = 12'h764;
        15'h1697: data = 12'h753;
        15'h1698: data = 12'h77A;
        15'h1699: data = 12'h7A3;
        15'h169A: data = 12'h7F1;
        15'h169B: data = 12'h0AA;
        15'h169C: data = 12'h10A;
        15'h169D: data = 12'h182;
        15'h169E: data = 12'h210;
        15'h169F: data = 12'h2B1;
        15'h16A0: data = 12'h363;
        15'h16A1: data = 12'h428;
        15'h16A2: data = 12'h4F9;
        15'h16A3: data = 12'h50D;
        15'h16A4: data = 12'h6D4;
        15'h16A5: data = 12'h7D1;
        15'h16A6: data = 12'h108;
        15'h16A7: data = 12'h215;
        15'h16A8: data = 12'h322;
        15'h16A9: data = 12'h43D;
        15'h16AA: data = 12'h551;
        15'h16AB: data = 12'h673;
        15'h16AC: data = 12'h792;
        15'h16AD: data = 12'h0F7;
        15'h16AE: data = 12'h211;
        15'h16AF: data = 12'h33B;
        15'h16B0: data = 12'h459;
        15'h16B1: data = 12'h569;
        15'h16B2: data = 12'h670;
        15'h16B3: data = 12'h76B;
        15'h16B4: data = 12'h491;
        15'h16B5: data = 12'h170;
        15'h16B6: data = 12'h23B;
        15'h16B7: data = 12'h2F7;
        15'h16B8: data = 12'h3AF;
        15'h16B9: data = 12'h453;
        15'h16BA: data = 12'h4EA;
        15'h16BB: data = 12'h562;
        15'h16BC: data = 12'h5DA;
        15'h16BD: data = 12'h61B;
        15'h16BE: data = 12'h659;
        15'h16BF: data = 12'h68D;
        15'h16C0: data = 12'h692;
        15'h16C1: data = 12'h68F;
        15'h16C2: data = 12'h50D;
        15'h16C3: data = 12'h632;
        15'h16C4: data = 12'h5E3;
        15'h16C5: data = 12'h590;
        15'h16C6: data = 12'h52B;
        15'h16C7: data = 12'h4A7;
        15'h16C8: data = 12'h412;
        15'h16C9: data = 12'h36D;
        15'h16CA: data = 12'h2B2;
        15'h16CB: data = 12'h1E4;
        15'h16CC: data = 12'h10B;
        15'h16CD: data = 12'h01E;
        15'h16CE: data = 12'h6E4;
        15'h16CF: data = 12'h5E7;
        15'h16D0: data = 12'h4D8;
        15'h16D1: data = 12'h3C2;
        15'h16D2: data = 12'h2AA;
        15'h16D3: data = 12'h18F;
        15'h16D4: data = 12'h079;
        15'h16D5: data = 12'h704;
        15'h16D6: data = 12'h5F0;
        15'h16D7: data = 12'h4D6;
        15'h16D8: data = 12'h3B6;
        15'h16D9: data = 12'h2A0;
        15'h16DA: data = 12'h188;
        15'h16DB: data = 12'h081;
        15'h16DC: data = 12'h746;
        15'h16DD: data = 12'h657;
        15'h16DE: data = 12'h567;
        15'h16DF: data = 12'h494;
        15'h16E0: data = 12'h3C9;
        15'h16E1: data = 12'h50D;
        15'h16E2: data = 12'h26C;
        15'h16E3: data = 12'h1D8;
        15'h16E4: data = 12'h144;
        15'h16E5: data = 12'h0E6;
        15'h16E6: data = 12'h08E;
        15'h16E7: data = 12'h032;
        15'h16E8: data = 12'h79F;
        15'h16E9: data = 12'h777;
        15'h16EA: data = 12'h754;
        15'h16EB: data = 12'h770;
        15'h16EC: data = 12'h795;
        15'h16ED: data = 12'h7D6;
        15'h16EE: data = 12'h2C6;
        15'h16EF: data = 12'h0E6;
        15'h16F0: data = 12'h156;
        15'h16F1: data = 12'h1DF;
        15'h16F2: data = 12'h279;
        15'h16F3: data = 12'h330;
        15'h16F4: data = 12'h3E9;
        15'h16F5: data = 12'h4B9;
        15'h16F6: data = 12'h592;
        15'h16F7: data = 12'h67E;
        15'h16F8: data = 12'h772;
        15'h16F9: data = 12'h0D0;
        15'h16FA: data = 12'h1AD;
        15'h16FB: data = 12'h2CE;
        15'h16FC: data = 12'h3DE;
        15'h16FD: data = 12'h500;
        15'h16FE: data = 12'h61B;
        15'h16FF: data = 12'h734;
        15'h1700: data = 12'h50D;
        15'h1701: data = 12'h1B8;
        15'h1702: data = 12'h2D1;
        15'h1703: data = 12'h3ED;
        15'h1704: data = 12'h4FF;
        15'h1705: data = 12'h613;
        15'h1706: data = 12'h716;
        15'h1707: data = 12'h809;
        15'h1708: data = 12'h12A;
        15'h1709: data = 12'h1FC;
        15'h170A: data = 12'h2C8;
        15'h170B: data = 12'h376;
        15'h170C: data = 12'h41E;
        15'h170D: data = 12'h4AF;
        15'h170E: data = 12'h539;
        15'h170F: data = 12'h5AB;
        15'h1710: data = 12'h5FC;
        15'h1711: data = 12'h654;
        15'h1712: data = 12'h674;
        15'h1713: data = 12'h695;
        15'h1714: data = 12'h695;
        15'h1715: data = 12'h66F;
        15'h1716: data = 12'h64E;
        15'h1717: data = 12'h606;
        15'h1718: data = 12'h5B2;
        15'h1719: data = 12'h54B;
        15'h171A: data = 12'h4CA;
        15'h171B: data = 12'h440;
        15'h171C: data = 12'h399;
        15'h171D: data = 12'h2ED;
        15'h171E: data = 12'h228;
        15'h171F: data = 12'h50D;
        15'h1720: data = 12'h071;
        15'h1721: data = 12'h73E;
        15'h1722: data = 12'h63E;
        15'h1723: data = 12'h536;
        15'h1724: data = 12'h41D;
        15'h1725: data = 12'h30A;
        15'h1726: data = 12'h1ED;
        15'h1727: data = 12'h0D3;
        15'h1728: data = 12'h76B;
        15'h1729: data = 12'h64D;
        15'h172A: data = 12'h531;
        15'h172B: data = 12'h419;
        15'h172C: data = 12'h2FC;
        15'h172D: data = 12'h1E4;
        15'h172E: data = 12'h0DD;
        15'h172F: data = 12'h786;
        15'h1730: data = 12'h6AA;
        15'h1731: data = 12'h5B9;
        15'h1732: data = 12'h4DE;
        15'h1733: data = 12'h40B;
        15'h1734: data = 12'h346;
        15'h1735: data = 12'h299;
        15'h1736: data = 12'h1FF;
        15'h1737: data = 12'h179;
        15'h1738: data = 12'h108;
        15'h1739: data = 12'h0A4;
        15'h173A: data = 12'h045;
        15'h173B: data = 12'h79F;
        15'h173C: data = 12'h77C;
        15'h173D: data = 12'h754;
        15'h173E: data = 12'h50D;
        15'h173F: data = 12'h778;
        15'h1740: data = 12'h7B5;
        15'h1741: data = 12'h7F8;
        15'h1742: data = 12'h0BF;
        15'h1743: data = 12'h12A;
        15'h1744: data = 12'h1B8;
        15'h1745: data = 12'h254;
        15'h1746: data = 12'h2FB;
        15'h1747: data = 12'h3B7;
        15'h1748: data = 12'h47F;
        15'h1749: data = 12'h548;
        15'h174A: data = 12'h62F;
        15'h174B: data = 12'h719;
        15'h174C: data = 12'h81A;
        15'h174D: data = 12'h157;
        15'h174E: data = 12'h268;
        15'h174F: data = 12'h384;
        15'h1750: data = 12'h4A6;
        15'h1751: data = 12'h5B9;
        15'h1752: data = 12'h6E1;
        15'h1753: data = 12'h7F1;
        15'h1754: data = 12'h157;
        15'h1755: data = 12'h274;
        15'h1756: data = 12'h38C;
        15'h1757: data = 12'h4AB;
        15'h1758: data = 12'h5B6;
        15'h1759: data = 12'h6C5;
        15'h175A: data = 12'h7B6;
        15'h175B: data = 12'h0E4;
        15'h175C: data = 12'h1C0;
        15'h175D: data = 12'h50D;
        15'h175E: data = 12'h341;
        15'h175F: data = 12'h3EF;
        15'h1760: data = 12'h487;
        15'h1761: data = 12'h510;
        15'h1762: data = 12'h580;
        15'h1763: data = 12'h5E7;
        15'h1764: data = 12'h635;
        15'h1765: data = 12'h675;
        15'h1766: data = 12'h691;
        15'h1767: data = 12'h696;
        15'h1768: data = 12'h694;
        15'h1769: data = 12'h66A;
        15'h176A: data = 12'h62C;
        15'h176B: data = 12'h5D4;
        15'h176C: data = 12'h564;
        15'h176D: data = 12'h4FB;
        15'h176E: data = 12'h46F;
        15'h176F: data = 12'h3D5;
        15'h1770: data = 12'h327;
        15'h1771: data = 12'h26E;
        15'h1772: data = 12'h19C;
        15'h1773: data = 12'h0C3;
        15'h1774: data = 12'h791;
        15'h1775: data = 12'h69E;
        15'h1776: data = 12'h595;
        15'h1777: data = 12'h48B;
        15'h1778: data = 12'h367;
        15'h1779: data = 12'h249;
        15'h177A: data = 12'h12E;
        15'h177B: data = 12'h093;
        15'h177C: data = 12'h50D;
        15'h177D: data = 12'h58A;
        15'h177E: data = 12'h475;
        15'h177F: data = 12'h35E;
        15'h1780: data = 12'h246;
        15'h1781: data = 12'h12B;
        15'h1782: data = 12'h02B;
        15'h1783: data = 12'h6F7;
        15'h1784: data = 12'h605;
        15'h1785: data = 12'h520;
        15'h1786: data = 12'h454;
        15'h1787: data = 12'h388;
        15'h1788: data = 12'h2D4;
        15'h1789: data = 12'h22D;
        15'h178A: data = 12'h19B;
        15'h178B: data = 12'h117;
        15'h178C: data = 12'h0C6;
        15'h178D: data = 12'h068;
        15'h178E: data = 12'h76A;
        15'h178F: data = 12'h784;
        15'h1790: data = 12'h771;
        15'h1791: data = 12'h757;
        15'h1792: data = 12'h773;
        15'h1793: data = 12'h797;
        15'h1794: data = 12'h7E1;
        15'h1795: data = 12'h099;
        15'h1796: data = 12'h107;
        15'h1797: data = 12'h180;
        15'h1798: data = 12'h21B;
        15'h1799: data = 12'h2BD;
        15'h179A: data = 12'h372;
        15'h179B: data = 12'h50D;
        15'h179C: data = 12'h500;
        15'h179D: data = 12'h5E0;
        15'h179E: data = 12'h6D3;
        15'h179F: data = 12'h7C9;
        15'h17A0: data = 12'h0FB;
        15'h17A1: data = 12'h205;
        15'h17A2: data = 12'h31A;
        15'h17A3: data = 12'h441;
        15'h17A4: data = 12'h556;
        15'h17A5: data = 12'h67A;
        15'h17A6: data = 12'h79D;
        15'h17A7: data = 12'h102;
        15'h17A8: data = 12'h219;
        15'h17A9: data = 12'h334;
        15'h17AA: data = 12'h44F;
        15'h17AB: data = 12'h559;
        15'h17AC: data = 12'h663;
        15'h17AD: data = 12'h762;
        15'h17AE: data = 12'h2B7;
        15'h17AF: data = 12'h178;
        15'h17B0: data = 12'h24E;
        15'h17B1: data = 12'h310;
        15'h17B2: data = 12'h3BA;
        15'h17B3: data = 12'h455;
        15'h17B4: data = 12'h4E4;
        15'h17B5: data = 12'h558;
        15'h17B6: data = 12'h5C9;
        15'h17B7: data = 12'h60C;
        15'h17B8: data = 12'h653;
        15'h17B9: data = 12'h68C;
        15'h17BA: data = 12'h50D;
        15'h17BB: data = 12'h697;
        15'h17BC: data = 12'h673;
        15'h17BD: data = 12'h639;
        15'h17BE: data = 12'h5ED;
        15'h17BF: data = 12'h58E;
        15'h17C0: data = 12'h529;
        15'h17C1: data = 12'h49B;
        15'h17C2: data = 12'h408;
        15'h17C3: data = 12'h360;
        15'h17C4: data = 12'h2A9;
        15'h17C5: data = 12'h1E5;
        15'h17C6: data = 12'h108;
        15'h17C7: data = 12'h048;
        15'h17C8: data = 12'h6EC;
        15'h17C9: data = 12'h5E9;
        15'h17CA: data = 12'h4D5;
        15'h17CB: data = 12'h3C8;
        15'h17CC: data = 12'h2A6;
        15'h17CD: data = 12'h18A;
        15'h17CE: data = 12'h075;
        15'h17CF: data = 12'h6FB;
        15'h17D0: data = 12'h5E3;
        15'h17D1: data = 12'h4D2;
        15'h17D2: data = 12'h3AF;
        15'h17D3: data = 12'h29F;
        15'h17D4: data = 12'h18C;
        15'h17D5: data = 12'h088;
        15'h17D6: data = 12'h74F;
        15'h17D7: data = 12'h65F;
        15'h17D8: data = 12'h56C;
        15'h17D9: data = 12'h50D;
        15'h17DA: data = 12'h3C7;
        15'h17DB: data = 12'h308;
        15'h17DC: data = 12'h25F;
        15'h17DD: data = 12'h1D1;
        15'h17DE: data = 12'h141;
        15'h17DF: data = 12'h0E7;
        15'h17E0: data = 12'h08A;
        15'h17E1: data = 12'h038;
        15'h17E2: data = 12'h7A7;
        15'h17E3: data = 12'h77F;
        15'h17E4: data = 12'h757;
        15'h17E5: data = 12'h772;
        15'h17E6: data = 12'h792;
        15'h17E7: data = 12'h7D4;
        15'h17E8: data = 12'h26C;
        15'h17E9: data = 12'h0DE;
        15'h17EA: data = 12'h155;
        15'h17EB: data = 12'h1DC;
        15'h17EC: data = 12'h27D;
        15'h17ED: data = 12'h335;
        15'h17EE: data = 12'h3F4;
        15'h17EF: data = 12'h4C2;
        15'h17F0: data = 12'h594;
        15'h17F1: data = 12'h684;
        15'h17F2: data = 12'h76F;
        15'h17F3: data = 12'h10F;
        15'h17F4: data = 12'h1A6;
        15'h17F5: data = 12'h2C6;
        15'h17F6: data = 12'h3E0;
        15'h17F7: data = 12'h503;
        15'h17F8: data = 12'h50D;
        15'h17F9: data = 12'h736;
        15'h17FA: data = 12'h509;
        15'h17FB: data = 12'h1BC;
        15'h17FC: data = 12'h2D1;
        15'h17FD: data = 12'h3ED;
        15'h17FE: data = 12'h4FE;
        15'h17FF: data = 12'h609;
        15'h1800: data = 12'h70D;
        15'h1801: data = 12'h803;
        15'h1802: data = 12'h128;
        15'h1803: data = 12'h1FE;
        15'h1804: data = 12'h2C8;
        15'h1805: data = 12'h37D;
        15'h1806: data = 12'h422;
        15'h1807: data = 12'h4B0;
        15'h1808: data = 12'h539;
        15'h1809: data = 12'h5A5;
        15'h180A: data = 12'h5F0;
        15'h180B: data = 12'h647;
        15'h180C: data = 12'h673;
        15'h180D: data = 12'h698;
        15'h180E: data = 12'h697;
        15'h180F: data = 12'h679;
        15'h1810: data = 12'h655;
        15'h1811: data = 12'h60E;
        15'h1812: data = 12'h5B7;
        15'h1813: data = 12'h546;
        15'h1814: data = 12'h4C7;
        15'h1815: data = 12'h43D;
        15'h1816: data = 12'h394;
        15'h1817: data = 12'h50D;
        15'h1818: data = 12'h225;
        15'h1819: data = 12'h14D;
        15'h181A: data = 12'h070;
        15'h181B: data = 12'h740;
        15'h181C: data = 12'h644;
        15'h181D: data = 12'h541;
        15'h181E: data = 12'h429;
        15'h181F: data = 12'h30E;
        15'h1820: data = 12'h1EB;
        15'h1821: data = 12'h0CC;
        15'h1822: data = 12'h762;
        15'h1823: data = 12'h63C;
        15'h1824: data = 12'h520;
        15'h1825: data = 12'h410;
        15'h1826: data = 12'h2F9;
        15'h1827: data = 12'h1E1;
        15'h1828: data = 12'h0DD;
        15'h1829: data = 12'h779;
        15'h182A: data = 12'h6AE;
        15'h182B: data = 12'h5C6;
        15'h182C: data = 12'h4E1;
        15'h182D: data = 12'h408;
        15'h182E: data = 12'h347;
        15'h182F: data = 12'h291;
        15'h1830: data = 12'h1F2;
        15'h1831: data = 12'h16C;
        15'h1832: data = 12'h103;
        15'h1833: data = 12'h0A0;
        15'h1834: data = 12'h04A;
        15'h1835: data = 12'h7A3;
        15'h1836: data = 12'h50D;
        15'h1837: data = 12'h761;
        15'h1838: data = 12'h779;
        15'h1839: data = 12'h77E;
        15'h183A: data = 12'h7B6;
        15'h183B: data = 12'h7F4;
        15'h183C: data = 12'h0B5;
        15'h183D: data = 12'h11D;
        15'h183E: data = 12'h1B1;
        15'h183F: data = 12'h253;
        15'h1840: data = 12'h2F8;
        15'h1841: data = 12'h3B4;
        15'h1842: data = 12'h482;
        15'h1843: data = 12'h54F;
        15'h1844: data = 12'h635;
        15'h1845: data = 12'h71E;
        15'h1846: data = 12'h81B;
        15'h1847: data = 12'h150;
        15'h1848: data = 12'h25F;
        15'h1849: data = 12'h37F;
        15'h184A: data = 12'h4A2;
        15'h184B: data = 12'h5B9;
        15'h184C: data = 12'h6E3;
        15'h184D: data = 12'h7FC;
        15'h184E: data = 12'h160;
        15'h184F: data = 12'h27F;
        15'h1850: data = 12'h393;
        15'h1851: data = 12'h4A7;
        15'h1852: data = 12'h5AD;
        15'h1853: data = 12'h6B8;
        15'h1854: data = 12'h7B1;
        15'h1855: data = 12'h50D;
        15'h1856: data = 12'h1BD;
        15'h1857: data = 12'h291;
        15'h1858: data = 12'h344;
        15'h1859: data = 12'h3FD;
        15'h185A: data = 12'h492;
        15'h185B: data = 12'h513;
        15'h185C: data = 12'h581;
        15'h185D: data = 12'h5E7;
        15'h185E: data = 12'h62A;
        15'h185F: data = 12'h671;
        15'h1860: data = 12'h694;
        15'h1861: data = 12'h697;
        15'h1862: data = 12'h695;
        15'h1863: data = 12'h672;
        15'h1864: data = 12'h638;
        15'h1865: data = 12'h5D7;
        15'h1866: data = 12'h56A;
        15'h1867: data = 12'h4FA;
        15'h1868: data = 12'h46D;
        15'h1869: data = 12'h3D2;
        15'h186A: data = 12'h326;
        15'h186B: data = 12'h264;
        15'h186C: data = 12'h19A;
        15'h186D: data = 12'h0BE;
        15'h186E: data = 12'h78D;
        15'h186F: data = 12'h699;
        15'h1870: data = 12'h591;
        15'h1871: data = 12'h486;
        15'h1872: data = 12'h364;
        15'h1873: data = 12'h24D;
        15'h1874: data = 12'h50D;
        15'h1875: data = 12'h039;
        15'h1876: data = 12'h69F;
        15'h1877: data = 12'h57E;
        15'h1878: data = 12'h46C;
        15'h1879: data = 12'h353;
        15'h187A: data = 12'h23D;
        15'h187B: data = 12'h12E;
        15'h187C: data = 12'h02D;
        15'h187D: data = 12'h6FF;
        15'h187E: data = 12'h60D;
        15'h187F: data = 12'h527;
        15'h1880: data = 12'h455;
        15'h1881: data = 12'h385;
        15'h1882: data = 12'h2D3;
        15'h1883: data = 12'h22A;
        15'h1884: data = 12'h194;
        15'h1885: data = 12'h114;
        15'h1886: data = 12'h0C2;
        15'h1887: data = 12'h067;
        15'h1888: data = 12'h759;
        15'h1889: data = 12'h783;
        15'h188A: data = 12'h771;
        15'h188B: data = 12'h75C;
        15'h188C: data = 12'h775;
        15'h188D: data = 12'h799;
        15'h188E: data = 12'h7E3;
        15'h188F: data = 12'h099;
        15'h1890: data = 12'h100;
        15'h1891: data = 12'h17A;
        15'h1892: data = 12'h20E;
        15'h1893: data = 12'h50D;
        15'h1894: data = 12'h371;
        15'h1895: data = 12'h439;
        15'h1896: data = 12'h50B;
        15'h1897: data = 12'h5E8;
        15'h1898: data = 12'h6D6;
        15'h1899: data = 12'h7C6;
        15'h189A: data = 12'h0FB;
        15'h189B: data = 12'h201;
        15'h189C: data = 12'h313;
        15'h189D: data = 12'h43A;
        15'h189E: data = 12'h553;
        15'h189F: data = 12'h67D;
        15'h18A0: data = 12'h79F;
        15'h18A1: data = 12'h109;
        15'h18A2: data = 12'h21D;
        15'h18A3: data = 12'h337;
        15'h18A4: data = 12'h449;
        15'h18A5: data = 12'h556;
        15'h18A6: data = 12'h65E;
        15'h18A7: data = 12'h75E;
        15'h18A8: data = 12'h1A6;
        15'h18A9: data = 12'h179;
        15'h18AA: data = 12'h24D;
        15'h18AB: data = 12'h30D;
        15'h18AC: data = 12'h3C6;
        15'h18AD: data = 12'h45F;
        15'h18AE: data = 12'h4EA;
        15'h18AF: data = 12'h55C;
        15'h18B0: data = 12'h5C5;
        15'h18B1: data = 12'h60A;
        15'h18B2: data = 12'h50D;
        15'h18B3: data = 12'h688;
        15'h18B4: data = 12'h694;
        15'h18B5: data = 12'h699;
        15'h18B6: data = 12'h675;
        15'h18B7: data = 12'h63C;
        15'h18B8: data = 12'h5F1;
        15'h18B9: data = 12'h595;
        15'h18BA: data = 12'h528;
        15'h18BB: data = 12'h49B;
        15'h18BC: data = 12'h404;
        15'h18BD: data = 12'h357;
        15'h18BE: data = 12'h2A1;
        15'h18BF: data = 12'h1DA;
        15'h18C0: data = 12'h105;
        15'h18C1: data = 12'h17B;
        15'h18C2: data = 12'h6ED;
        15'h18C3: data = 12'h5F1;
        15'h18C4: data = 12'h4E3;
        15'h18C5: data = 12'h3CE;
        15'h18C6: data = 12'h2AE;
        15'h18C7: data = 12'h18D;
        15'h18C8: data = 12'h06E;
        15'h18C9: data = 12'h6F7;
        15'h18CA: data = 12'h5E4;
        15'h18CB: data = 12'h4CE;
        15'h18CC: data = 12'h3AA;
        15'h18CD: data = 12'h29F;
        15'h18CE: data = 12'h187;
        15'h18CF: data = 12'h086;
        15'h18D0: data = 12'h74F;
        15'h18D1: data = 12'h50D;
        15'h18D2: data = 12'h56E;
        15'h18D3: data = 12'h497;
        15'h18D4: data = 12'h3CA;
        15'h18D5: data = 12'h309;
        15'h18D6: data = 12'h25F;
        15'h18D7: data = 12'h1C8;
        15'h18D8: data = 12'h136;
        15'h18D9: data = 12'h0E1;
        15'h18DA: data = 12'h085;
        15'h18DB: data = 12'h037;
        15'h18DC: data = 12'h7A8;
        15'h18DD: data = 12'h783;
        15'h18DE: data = 12'h760;
        15'h18DF: data = 12'h779;
        15'h18E0: data = 12'h793;
        15'h18E1: data = 12'h7D3;
        15'h18E2: data = 12'h290;
        15'h18E3: data = 12'h0DB;
        15'h18E4: data = 12'h14F;
        15'h18E5: data = 12'h1DF;
        15'h18E6: data = 12'h27F;
        15'h18E7: data = 12'h337;
        15'h18E8: data = 12'h3F5;
        15'h18E9: data = 12'h4C3;
        15'h18EA: data = 12'h59F;
        15'h18EB: data = 12'h688;
        15'h18EC: data = 12'h774;
        15'h18ED: data = 12'h10A;
        15'h18EE: data = 12'h1A2;
        15'h18EF: data = 12'h2C1;
        15'h18F0: data = 12'h50D;
        15'h18F1: data = 12'h504;
        15'h18F2: data = 12'h621;
        15'h18F3: data = 12'h737;
        15'h18F4: data = 12'h556;
        15'h18F5: data = 12'h1C7;
        15'h18F6: data = 12'h2D7;
        15'h18F7: data = 12'h3F3;
        15'h18F8: data = 12'h502;
        15'h18F9: data = 12'h60A;
        15'h18FA: data = 12'h710;
        15'h18FB: data = 12'h807;
        15'h18FC: data = 12'h129;
        15'h18FD: data = 12'h204;
        15'h18FE: data = 12'h2D1;
        15'h18FF: data = 12'h385;
        15'h1900: data = 12'h42E;
        15'h1901: data = 12'h4BB;
        15'h1902: data = 12'h543;
        15'h1903: data = 12'h5A0;
        15'h1904: data = 12'h5F2;
        15'h1905: data = 12'h647;
        15'h1906: data = 12'h66D;
        15'h1907: data = 12'h695;
        15'h1908: data = 12'h695;
        15'h1909: data = 12'h679;
        15'h190A: data = 12'h659;
        15'h190B: data = 12'h614;
        15'h190C: data = 12'h5BB;
        15'h190D: data = 12'h54D;
        15'h190E: data = 12'h4C8;
        15'h190F: data = 12'h50D;
        15'h1910: data = 12'h393;
        15'h1911: data = 12'h2E1;
        15'h1912: data = 12'h21C;
        15'h1913: data = 12'h148;
        15'h1914: data = 12'h071;
        15'h1915: data = 12'h740;
        15'h1916: data = 12'h642;
        15'h1917: data = 12'h53B;
        15'h1918: data = 12'h427;
        15'h1919: data = 12'h318;
        15'h191A: data = 12'h1F3;
        15'h191B: data = 12'h0CF;
        15'h191C: data = 12'h767;
        15'h191D: data = 12'h63B;
        15'h191E: data = 12'h51A;
        15'h191F: data = 12'h40A;
        15'h1920: data = 12'h2FA;
        15'h1921: data = 12'h1E3;
        15'h1922: data = 12'h0DB;
        15'h1923: data = 12'h765;
        15'h1924: data = 12'h6B4;
        15'h1925: data = 12'h5C2;
        15'h1926: data = 12'h4E5;
        15'h1927: data = 12'h40C;
        15'h1928: data = 12'h347;
        15'h1929: data = 12'h291;
        15'h192A: data = 12'h1F2;
        15'h192B: data = 12'h16A;
        15'h192C: data = 12'h0FB;
        15'h192D: data = 12'h099;
        15'h192E: data = 12'h50D;
        15'h192F: data = 12'h7A2;
        15'h1930: data = 12'h787;
        15'h1931: data = 12'h761;
        15'h1932: data = 12'h784;
        15'h1933: data = 12'h784;
        15'h1934: data = 12'h7B4;
        15'h1935: data = 12'h7F5;
        15'h1936: data = 12'h0B4;
        15'h1937: data = 12'h11E;
        15'h1938: data = 12'h1AD;
        15'h1939: data = 12'h24D;
        15'h193A: data = 12'h2F9;
        15'h193B: data = 12'h3B8;
        15'h193C: data = 12'h486;
        15'h193D: data = 12'h54F;
        15'h193E: data = 12'h638;
        15'h193F: data = 12'h722;
        15'h1940: data = 12'h81A;
        15'h1941: data = 12'h14F;
        15'h1942: data = 12'h260;
        15'h1943: data = 12'h378;
        15'h1944: data = 12'h499;
        15'h1945: data = 12'h5B3;
        15'h1946: data = 12'h6E0;
        15'h1947: data = 12'h7FD;
        15'h1948: data = 12'h167;
        15'h1949: data = 12'h28A;
        15'h194A: data = 12'h399;
        15'h194B: data = 12'h4AB;
        15'h194C: data = 12'h5AC;
        15'h194D: data = 12'h50D;
        15'h194E: data = 12'h7A5;
        15'h194F: data = 12'h0D9;
        15'h1950: data = 12'h1B7;
        15'h1951: data = 12'h291;
        15'h1952: data = 12'h346;
        15'h1953: data = 12'h3FB;
        15'h1954: data = 12'h496;
        15'h1955: data = 12'h519;
        15'h1956: data = 12'h585;
        15'h1957: data = 12'h5E8;
        15'h1958: data = 12'h629;
        15'h1959: data = 12'h667;
        15'h195A: data = 12'h688;
        15'h195B: data = 12'h68D;
        15'h195C: data = 12'h693;
        15'h195D: data = 12'h673;
        15'h195E: data = 12'h636;
        15'h195F: data = 12'h5DB;
        15'h1960: data = 12'h571;
        15'h1961: data = 12'h502;
        15'h1962: data = 12'h472;
        15'h1963: data = 12'h3D2;
        15'h1964: data = 12'h31C;
        15'h1965: data = 12'h25B;
        15'h1966: data = 12'h18C;
        15'h1967: data = 12'h0AF;
        15'h1968: data = 12'h788;
        15'h1969: data = 12'h697;
        15'h196A: data = 12'h590;
        15'h196B: data = 12'h48A;
        15'h196C: data = 12'h50D;
        15'h196D: data = 12'h258;
        15'h196E: data = 12'h137;
        15'h196F: data = 12'h015;
        15'h1970: data = 12'h6A1;
        15'h1971: data = 12'h579;
        15'h1972: data = 12'h464;
        15'h1973: data = 12'h348;
        15'h1974: data = 12'h234;
        15'h1975: data = 12'h126;
        15'h1976: data = 12'h093;
        15'h1977: data = 12'h700;
        15'h1978: data = 12'h610;
        15'h1979: data = 12'h533;
        15'h197A: data = 12'h465;
        15'h197B: data = 12'h393;
        15'h197C: data = 12'h2D4;
        15'h197D: data = 12'h22B;
        15'h197E: data = 12'h18E;
        15'h197F: data = 12'h108;
        15'h1980: data = 12'h0B2;
        15'h1981: data = 12'h059;
        15'h1982: data = 12'h7C3;
        15'h1983: data = 12'h782;
        15'h1984: data = 12'h778;
        15'h1985: data = 12'h766;
        15'h1986: data = 12'h782;
        15'h1987: data = 12'h7A6;
        15'h1988: data = 12'h7EC;
        15'h1989: data = 12'h094;
        15'h198A: data = 12'h0FD;
        15'h198B: data = 12'h50D;
        15'h198C: data = 12'h204;
        15'h198D: data = 12'h2AB;
        15'h198E: data = 12'h368;
        15'h198F: data = 12'h438;
        15'h1990: data = 12'h50B;
        15'h1991: data = 12'h5F1;
        15'h1992: data = 12'h6E0;
        15'h1993: data = 12'h7D7;
        15'h1994: data = 12'h104;
        15'h1995: data = 12'h208;
        15'h1996: data = 12'h30D;
        15'h1997: data = 12'h430;
        15'h1998: data = 12'h54A;
        15'h1999: data = 12'h675;
        15'h199A: data = 12'h79D;
        15'h199B: data = 12'h10D;
        15'h199C: data = 12'h222;
        15'h199D: data = 12'h343;
        15'h199E: data = 12'h455;
        15'h199F: data = 12'h560;
        15'h19A0: data = 12'h65F;
        15'h19A1: data = 12'h759;
        15'h19A2: data = 12'h20F;
        15'h19A3: data = 12'h165;
        15'h19A4: data = 12'h23F;
        15'h19A5: data = 12'h307;
        15'h19A6: data = 12'h3C0;
        15'h19A7: data = 12'h464;
        15'h19A8: data = 12'h4F5;
        15'h19A9: data = 12'h56B;
        15'h19AA: data = 12'h50D;
        15'h19AB: data = 12'h60F;
        15'h19AC: data = 12'h646;
        15'h19AD: data = 12'h67D;
        15'h19AE: data = 12'h683;
        15'h19AF: data = 12'h687;
        15'h19B0: data = 12'h66D;
        15'h19B1: data = 12'h63D;
        15'h19B2: data = 12'h5F4;
        15'h19B3: data = 12'h59A;
        15'h19B4: data = 12'h535;
        15'h19B5: data = 12'h4A6;
        15'h19B6: data = 12'h40B;
        15'h19B7: data = 12'h35C;
        15'h19B8: data = 12'h2A2;
        15'h19B9: data = 12'h1D5;
        15'h19BA: data = 12'h0FA;
        15'h19BB: data = 12'h08F;
        15'h19BC: data = 12'h6E5;
        15'h19BD: data = 12'h5EA;
        15'h19BE: data = 12'h4DF;
        15'h19BF: data = 12'h3D0;
        15'h19C0: data = 12'h2B5;
        15'h19C1: data = 12'h197;
        15'h19C2: data = 12'h07D;
        15'h19C3: data = 12'h702;
        15'h19C4: data = 12'h5E4;
        15'h19C5: data = 12'h4C9;
        15'h19C6: data = 12'h3A0;
        15'h19C7: data = 12'h28A;
        15'h19C8: data = 12'h172;
        15'h19C9: data = 12'h50D;
        15'h19CA: data = 12'h74A;
        15'h19CB: data = 12'h667;
        15'h19CC: data = 12'h576;
        15'h19CD: data = 12'h4A8;
        15'h19CE: data = 12'h3D7;
        15'h19CF: data = 12'h31C;
        15'h19D0: data = 12'h26A;
        15'h19D1: data = 12'h1D1;
        15'h19D2: data = 12'h137;
        15'h19D3: data = 12'h0D5;
        15'h19D4: data = 12'h078;
        15'h19D5: data = 12'h025;
        15'h19D6: data = 12'h799;
        15'h19D7: data = 12'h77F;
        15'h19D8: data = 12'h763;
        15'h19D9: data = 12'h786;
        15'h19DA: data = 12'h7A6;
        15'h19DB: data = 12'h7E3;
        15'h19DC: data = 12'h737;
        15'h19DD: data = 12'h0DF;
        15'h19DE: data = 12'h14A;
        15'h19DF: data = 12'h1CF;
        15'h19E0: data = 12'h26F;
        15'h19E1: data = 12'h329;
        15'h19E2: data = 12'h3ED;
        15'h19E3: data = 12'h4C3;
        15'h19E4: data = 12'h59F;
        15'h19E5: data = 12'h68E;
        15'h19E6: data = 12'h77F;
        15'h19E7: data = 12'h0AB;
        15'h19E8: data = 12'h50D;
        15'h19E9: data = 12'h2C2;
        15'h19EA: data = 12'h3D5;
        15'h19EB: data = 12'h4F8;
        15'h19EC: data = 12'h613;
        15'h19ED: data = 12'h72D;
        15'h19EE: data = 12'h277;
        15'h19EF: data = 12'h1C1;
        15'h19F0: data = 12'h2E5;
        15'h19F1: data = 12'h401;
        15'h19F2: data = 12'h513;
        15'h19F3: data = 12'h619;
        15'h19F4: data = 12'h714;
        15'h19F5: data = 12'h7FC;
        15'h19F6: data = 12'h119;
        15'h19F7: data = 12'h1EE;
        15'h19F8: data = 12'h2C1;
        15'h19F9: data = 12'h37C;
        15'h19FA: data = 12'h42B;
        15'h19FB: data = 12'h4C4;
        15'h19FC: data = 12'h550;
        15'h19FD: data = 12'h5B9;
        15'h19FE: data = 12'h603;
        15'h19FF: data = 12'h64E;
        15'h1A00: data = 12'h66A;
        15'h1A01: data = 12'h686;
        15'h1A02: data = 12'h688;
        15'h1A03: data = 12'h663;
        15'h1A04: data = 12'h649;
        15'h1A05: data = 12'h610;
        15'h1A06: data = 12'h5BF;
        15'h1A07: data = 12'h50D;
        15'h1A08: data = 12'h4E3;
        15'h1A09: data = 12'h44A;
        15'h1A0A: data = 12'h3A4;
        15'h1A0B: data = 12'h2EA;
        15'h1A0C: data = 12'h21A;
        15'h1A0D: data = 12'h13E;
        15'h1A0E: data = 12'h05F;
        15'h1A0F: data = 12'h729;
        15'h1A10: data = 12'h631;
        15'h1A11: data = 12'h52F;
        15'h1A12: data = 12'h424;
        15'h1A13: data = 12'h318;
        15'h1A14: data = 12'h1FF;
        15'h1A15: data = 12'h0DC;
        15'h1A16: data = 12'h771;
        15'h1A17: data = 12'h64A;
        15'h1A18: data = 12'h525;
        15'h1A19: data = 12'h409;
        15'h1A1A: data = 12'h2E6;
        15'h1A1B: data = 12'h1D0;
        15'h1A1C: data = 12'h0C9;
        15'h1A1D: data = 12'h79E;
        15'h1A1E: data = 12'h6A8;
        15'h1A1F: data = 12'h5BE;
        15'h1A20: data = 12'h4E4;
        15'h1A21: data = 12'h414;
        15'h1A22: data = 12'h357;
        15'h1A23: data = 12'h2A3;
        15'h1A24: data = 12'h1FF;
        15'h1A25: data = 12'h178;
        15'h1A26: data = 12'h50D;
        15'h1A27: data = 12'h091;
        15'h1A28: data = 12'h037;
        15'h1A29: data = 12'h793;
        15'h1A2A: data = 12'h772;
        15'h1A2B: data = 12'h753;
        15'h1A2C: data = 12'h77C;
        15'h1A2D: data = 12'h783;
        15'h1A2E: data = 12'h7C3;
        15'h1A2F: data = 12'h807;
        15'h1A30: data = 12'h0C6;
        15'h1A31: data = 12'h131;
        15'h1A32: data = 12'h1B6;
        15'h1A33: data = 12'h246;
        15'h1A34: data = 12'h2E9;
        15'h1A35: data = 12'h3A0;
        15'h1A36: data = 12'h471;
        15'h1A37: data = 12'h542;
        15'h1A38: data = 12'h637;
        15'h1A39: data = 12'h72C;
        15'h1A3A: data = 12'h82C;
        15'h1A3B: data = 12'h164;
        15'h1A3C: data = 12'h270;
        15'h1A3D: data = 12'h386;
        15'h1A3E: data = 12'h49A;
        15'h1A3F: data = 12'h5AB;
        15'h1A40: data = 12'h6D2;
        15'h1A41: data = 12'h7E9;
        15'h1A42: data = 12'h157;
        15'h1A43: data = 12'h27D;
        15'h1A44: data = 12'h39D;
        15'h1A45: data = 12'h50D;
        15'h1A46: data = 12'h5C0;
        15'h1A47: data = 12'h6C7;
        15'h1A48: data = 12'h7B9;
        15'h1A49: data = 12'h0E1;
        15'h1A4A: data = 12'h1B3;
        15'h1A4B: data = 12'h285;
        15'h1A4C: data = 12'h339;
        15'h1A4D: data = 12'h3ED;
        15'h1A4E: data = 12'h490;
        15'h1A4F: data = 12'h519;
        15'h1A50: data = 12'h58F;
        15'h1A51: data = 12'h5FC;
        15'h1A52: data = 12'h63C;
        15'h1A53: data = 12'h679;
        15'h1A54: data = 12'h695;
        15'h1A55: data = 12'h691;
        15'h1A56: data = 12'h688;
        15'h1A57: data = 12'h65E;
        15'h1A58: data = 12'h628;
        15'h1A59: data = 12'h5D2;
        15'h1A5A: data = 12'h56C;
        15'h1A5B: data = 12'h4FF;
        15'h1A5C: data = 12'h47D;
        15'h1A5D: data = 12'h3E5;
        15'h1A5E: data = 12'h336;
        15'h1A5F: data = 12'h26C;
        15'h1A60: data = 12'h199;
        15'h1A61: data = 12'h0B4;
        15'h1A62: data = 12'h787;
        15'h1A63: data = 12'h689;
        15'h1A64: data = 12'h50D;
        15'h1A65: data = 12'h47E;
        15'h1A66: data = 12'h364;
        15'h1A67: data = 12'h24F;
        15'h1A68: data = 12'h138;
        15'h1A69: data = 12'h210;
        15'h1A6A: data = 12'h6B1;
        15'h1A6B: data = 12'h58A;
        15'h1A6C: data = 12'h474;
        15'h1A6D: data = 12'h34F;
        15'h1A6E: data = 12'h23B;
        15'h1A6F: data = 12'h123;
        15'h1A70: data = 12'h01F;
        15'h1A71: data = 12'h6ED;
        15'h1A72: data = 12'h5FD;
        15'h1A73: data = 12'h521;
        15'h1A74: data = 12'h453;
        15'h1A75: data = 12'h38A;
        15'h1A76: data = 12'h2DE;
        15'h1A77: data = 12'h23C;
        15'h1A78: data = 12'h1A6;
        15'h1A79: data = 12'h11F;
        15'h1A7A: data = 12'h0C0;
        15'h1A7B: data = 12'h060;
        15'h1A7C: data = 12'h7A2;
        15'h1A7D: data = 12'h773;
        15'h1A7E: data = 12'h763;
        15'h1A7F: data = 12'h751;
        15'h1A80: data = 12'h776;
        15'h1A81: data = 12'h7A2;
        15'h1A82: data = 12'h7EF;
        15'h1A83: data = 12'h50D;
        15'h1A84: data = 12'h111;
        15'h1A85: data = 12'h181;
        15'h1A86: data = 12'h213;
        15'h1A87: data = 12'h2B5;
        15'h1A88: data = 12'h366;
        15'h1A89: data = 12'h428;
        15'h1A8A: data = 12'h4FB;
        15'h1A8B: data = 12'h5E2;
        15'h1A8C: data = 12'h6D6;
        15'h1A8D: data = 12'h7D5;
        15'h1A8E: data = 12'h10A;
        15'h1A8F: data = 12'h218;
        15'h1A90: data = 12'h321;
        15'h1A91: data = 12'h440;
        15'h1A92: data = 12'h556;
        15'h1A93: data = 12'h675;
        15'h1A94: data = 12'h793;
        15'h1A95: data = 12'h101;
        15'h1A96: data = 12'h217;
        15'h1A97: data = 12'h338;
        15'h1A98: data = 12'h453;
        15'h1A99: data = 12'h564;
        15'h1A9A: data = 12'h66F;
        15'h1A9B: data = 12'h76B;
        15'h1A9C: data = 12'h457;
        15'h1A9D: data = 12'h17B;
        15'h1A9E: data = 12'h248;
        15'h1A9F: data = 12'h304;
        15'h1AA0: data = 12'h3B2;
        15'h1AA1: data = 12'h44E;
        15'h1AA2: data = 12'h50D;
        15'h1AA3: data = 12'h560;
        15'h1AA4: data = 12'h5D2;
        15'h1AA5: data = 12'h619;
        15'h1AA6: data = 12'h658;
        15'h1AA7: data = 12'h690;
        15'h1AA8: data = 12'h696;
        15'h1AA9: data = 12'h690;
        15'h1AAA: data = 12'h66A;
        15'h1AAB: data = 12'h631;
        15'h1AAC: data = 12'h5E7;
        15'h1AAD: data = 12'h58E;
        15'h1AAE: data = 12'h52D;
        15'h1AAF: data = 12'h49F;
        15'h1AB0: data = 12'h40F;
        15'h1AB1: data = 12'h365;
        15'h1AB2: data = 12'h2AD;
        15'h1AB3: data = 12'h1E4;
        15'h1AB4: data = 12'h10A;
        15'h1AB5: data = 12'h01F;
        15'h1AB6: data = 12'h6E3;
        15'h1AB7: data = 12'h5E1;
        15'h1AB8: data = 12'h4D3;
        15'h1AB9: data = 12'h3BD;
        15'h1ABA: data = 12'h2A4;
        15'h1ABB: data = 12'h18E;
        15'h1ABC: data = 12'h074;
        15'h1ABD: data = 12'h704;
        15'h1ABE: data = 12'h5F0;
        15'h1ABF: data = 12'h4D9;
        15'h1AC0: data = 12'h3B3;
        15'h1AC1: data = 12'h50D;
        15'h1AC2: data = 12'h186;
        15'h1AC3: data = 12'h07F;
        15'h1AC4: data = 12'h741;
        15'h1AC5: data = 12'h655;
        15'h1AC6: data = 12'h560;
        15'h1AC7: data = 12'h491;
        15'h1AC8: data = 12'h3C5;
        15'h1AC9: data = 12'h30F;
        15'h1ACA: data = 12'h26A;
        15'h1ACB: data = 12'h1D2;
        15'h1ACC: data = 12'h141;
        15'h1ACD: data = 12'h0E9;
        15'h1ACE: data = 12'h08A;
        15'h1ACF: data = 12'h02E;
        15'h1AD0: data = 12'h79A;
        15'h1AD1: data = 12'h776;
        15'h1AD2: data = 12'h753;
        15'h1AD3: data = 12'h770;
        15'h1AD4: data = 12'h794;
        15'h1AD5: data = 12'h7D4;
        15'h1AD6: data = 12'h22D;
        15'h1AD7: data = 12'h0E4;
        15'h1AD8: data = 12'h15C;
        15'h1AD9: data = 12'h1E3;
        15'h1ADA: data = 12'h27F;
        15'h1ADB: data = 12'h336;
        15'h1ADC: data = 12'h3F6;
        15'h1ADD: data = 12'h4C1;
        15'h1ADE: data = 12'h593;
        15'h1ADF: data = 12'h67E;
        15'h1AE0: data = 12'h50D;
        15'h1AE1: data = 12'h0E2;
        15'h1AE2: data = 12'h1AB;
        15'h1AE3: data = 12'h2CF;
        15'h1AE4: data = 12'h3E8;
        15'h1AE5: data = 12'h507;
        15'h1AE6: data = 12'h622;
        15'h1AE7: data = 12'h735;
        15'h1AE8: data = 12'h437;
        15'h1AE9: data = 12'h1BC;
        15'h1AEA: data = 12'h2D7;
        15'h1AEB: data = 12'h3F0;
        15'h1AEC: data = 12'h509;
        15'h1AED: data = 12'h611;
        15'h1AEE: data = 12'h714;
        15'h1AEF: data = 12'h80D;
        15'h1AF0: data = 12'h131;
        15'h1AF1: data = 12'h203;
        15'h1AF2: data = 12'h2D0;
        15'h1AF3: data = 12'h37E;
        15'h1AF4: data = 12'h424;
        15'h1AF5: data = 12'h4B3;
        15'h1AF6: data = 12'h53D;
        15'h1AF7: data = 12'h5A6;
        15'h1AF8: data = 12'h5FC;
        15'h1AF9: data = 12'h64F;
        15'h1AFA: data = 12'h676;
        15'h1AFB: data = 12'h697;
        15'h1AFC: data = 12'h697;
        15'h1AFD: data = 12'h678;
        15'h1AFE: data = 12'h655;
        15'h1AFF: data = 12'h50D;
        15'h1B00: data = 12'h5B3;
        15'h1B01: data = 12'h549;
        15'h1B02: data = 12'h4CB;
        15'h1B03: data = 12'h43B;
        15'h1B04: data = 12'h39A;
        15'h1B05: data = 12'h2EC;
        15'h1B06: data = 12'h228;
        15'h1B07: data = 12'h150;
        15'h1B08: data = 12'h073;
        15'h1B09: data = 12'h740;
        15'h1B0A: data = 12'h640;
        15'h1B0B: data = 12'h539;
        15'h1B0C: data = 12'h41D;
        15'h1B0D: data = 12'h30C;
        15'h1B0E: data = 12'h1EB;
        15'h1B0F: data = 12'h0CD;
        15'h1B10: data = 12'h763;
        15'h1B11: data = 12'h63F;
        15'h1B12: data = 12'h521;
        15'h1B13: data = 12'h412;
        15'h1B14: data = 12'h2FB;
        15'h1B15: data = 12'h1E3;
        15'h1B16: data = 12'h0E0;
        15'h1B17: data = 12'h787;
        15'h1B18: data = 12'h6AC;
        15'h1B19: data = 12'h5B9;
        15'h1B1A: data = 12'h4E0;
        15'h1B1B: data = 12'h40A;
        15'h1B1C: data = 12'h347;
        15'h1B1D: data = 12'h292;
        15'h1B1E: data = 12'h50D;
        15'h1B1F: data = 12'h172;
        15'h1B20: data = 12'h105;
        15'h1B21: data = 12'h0A3;
        15'h1B22: data = 12'h046;
        15'h1B23: data = 12'h7A2;
        15'h1B24: data = 12'h784;
        15'h1B25: data = 12'h75B;
        15'h1B26: data = 12'h777;
        15'h1B27: data = 12'h778;
        15'h1B28: data = 12'h7B3;
        15'h1B29: data = 12'h7F9;
        15'h1B2A: data = 12'h0B5;
        15'h1B2B: data = 12'h12A;
        15'h1B2C: data = 12'h1B9;
        15'h1B2D: data = 12'h254;
        15'h1B2E: data = 12'h2FE;
        15'h1B2F: data = 12'h3B3;
        15'h1B30: data = 12'h481;
        15'h1B31: data = 12'h549;
        15'h1B32: data = 12'h630;
        15'h1B33: data = 12'h719;
        15'h1B34: data = 12'h818;
        15'h1B35: data = 12'h14E;
        15'h1B36: data = 12'h26B;
        15'h1B37: data = 12'h387;
        15'h1B38: data = 12'h4A7;
        15'h1B39: data = 12'h5BD;
        15'h1B3A: data = 12'h6E6;
        15'h1B3B: data = 12'h7F7;
        15'h1B3C: data = 12'h15E;
        15'h1B3D: data = 12'h50D;
        15'h1B3E: data = 12'h38B;
        15'h1B3F: data = 12'h4A6;
        15'h1B40: data = 12'h5B2;
        15'h1B41: data = 12'h6BC;
        15'h1B42: data = 12'h7B0;
        15'h1B43: data = 12'h0E5;
        15'h1B44: data = 12'h1BF;
        15'h1B45: data = 12'h28F;
        15'h1B46: data = 12'h346;
        15'h1B47: data = 12'h3F5;
        15'h1B48: data = 12'h490;
        15'h1B49: data = 12'h512;
        15'h1B4A: data = 12'h57F;
        15'h1B4B: data = 12'h5E8;
        15'h1B4C: data = 12'h627;
        15'h1B4D: data = 12'h670;
        15'h1B4E: data = 12'h699;
        15'h1B4F: data = 12'h699;
        15'h1B50: data = 12'h698;
        15'h1B51: data = 12'h66E;
        15'h1B52: data = 12'h631;
        15'h1B53: data = 12'h5D3;
        15'h1B54: data = 12'h567;
        15'h1B55: data = 12'h4F4;
        15'h1B56: data = 12'h46E;
        15'h1B57: data = 12'h3D1;
        15'h1B58: data = 12'h328;
        15'h1B59: data = 12'h26F;
        15'h1B5A: data = 12'h19D;
        15'h1B5B: data = 12'h0BF;
        15'h1B5C: data = 12'h50D;
        15'h1B5D: data = 12'h697;
        15'h1B5E: data = 12'h58D;
        15'h1B5F: data = 12'h484;
        15'h1B60: data = 12'h361;
        15'h1B61: data = 12'h247;
        15'h1B62: data = 12'h12E;
        15'h1B63: data = 12'h04E;
        15'h1B64: data = 12'h6A5;
        15'h1B65: data = 12'h585;
        15'h1B66: data = 12'h46F;
        15'h1B67: data = 12'h352;
        15'h1B68: data = 12'h23F;
        15'h1B69: data = 12'h12F;
        15'h1B6A: data = 12'h02C;
        15'h1B6B: data = 12'h6FF;
        15'h1B6C: data = 12'h60C;
        15'h1B6D: data = 12'h52A;
        15'h1B6E: data = 12'h456;
        15'h1B6F: data = 12'h385;
        15'h1B70: data = 12'h2D0;
        15'h1B71: data = 12'h228;
        15'h1B72: data = 12'h194;
        15'h1B73: data = 12'h114;
        15'h1B74: data = 12'h0C0;
        15'h1B75: data = 12'h069;
        15'h1B76: data = 12'h77E;
        15'h1B77: data = 12'h781;
        15'h1B78: data = 12'h772;
        15'h1B79: data = 12'h75C;
        15'h1B7A: data = 12'h778;
        15'h1B7B: data = 12'h50D;
        15'h1B7C: data = 12'h7E2;
        15'h1B7D: data = 12'h098;
        15'h1B7E: data = 12'h103;
        15'h1B7F: data = 12'h17D;
        15'h1B80: data = 12'h211;
        15'h1B81: data = 12'h2BD;
        15'h1B82: data = 12'h376;
        15'h1B83: data = 12'h43B;
        15'h1B84: data = 12'h509;
        15'h1B85: data = 12'h5E3;
        15'h1B86: data = 12'h6D1;
        15'h1B87: data = 12'h7C5;
        15'h1B88: data = 12'h0F7;
        15'h1B89: data = 12'h206;
        15'h1B8A: data = 12'h31B;
        15'h1B8B: data = 12'h443;
        15'h1B8C: data = 12'h55B;
        15'h1B8D: data = 12'h682;
        15'h1B8E: data = 12'h79E;
        15'h1B8F: data = 12'h106;
        15'h1B90: data = 12'h216;
        15'h1B91: data = 12'h332;
        15'h1B92: data = 12'h448;
        15'h1B93: data = 12'h556;
        15'h1B94: data = 12'h663;
        15'h1B95: data = 12'h766;
        15'h1B96: data = 12'h10D;
        15'h1B97: data = 12'h17A;
        15'h1B98: data = 12'h24C;
        15'h1B99: data = 12'h308;
        15'h1B9A: data = 12'h50D;
        15'h1B9B: data = 12'h456;
        15'h1B9C: data = 12'h4E5;
        15'h1B9D: data = 12'h559;
        15'h1B9E: data = 12'h5CA;
        15'h1B9F: data = 12'h60C;
        15'h1BA0: data = 12'h64C;
        15'h1BA1: data = 12'h689;
        15'h1BA2: data = 12'h698;
        15'h1BA3: data = 12'h69B;
        15'h1BA4: data = 12'h679;
        15'h1BA5: data = 12'h63D;
        15'h1BA6: data = 12'h5ED;
        15'h1BA7: data = 12'h592;
        15'h1BA8: data = 12'h52A;
        15'h1BA9: data = 12'h49C;
        15'h1BAA: data = 12'h409;
        15'h1BAB: data = 12'h35D;
        15'h1BAC: data = 12'h2A6;
        15'h1BAD: data = 12'h1DC;
        15'h1BAE: data = 12'h102;
        15'h1BAF: data = 12'h27F;
        15'h1BB0: data = 12'h6ED;
        15'h1BB1: data = 12'h5EB;
        15'h1BB2: data = 12'h4DE;
        15'h1BB3: data = 12'h3CA;
        15'h1BB4: data = 12'h2A9;
        15'h1BB5: data = 12'h187;
        15'h1BB6: data = 12'h06C;
        15'h1BB7: data = 12'h6FA;
        15'h1BB8: data = 12'h5E1;
        15'h1BB9: data = 12'h50D;
        15'h1BBA: data = 12'h3AD;
        15'h1BBB: data = 12'h2A3;
        15'h1BBC: data = 12'h18E;
        15'h1BBD: data = 12'h085;
        15'h1BBE: data = 12'h747;
        15'h1BBF: data = 12'h65D;
        15'h1BC0: data = 12'h56B;
        15'h1BC1: data = 12'h493;
        15'h1BC2: data = 12'h3C9;
        15'h1BC3: data = 12'h30B;
        15'h1BC4: data = 12'h260;
        15'h1BC5: data = 12'h1CB;
        15'h1BC6: data = 12'h13B;
        15'h1BC7: data = 12'h0E1;
        15'h1BC8: data = 12'h087;
        15'h1BC9: data = 12'h034;
        15'h1BCA: data = 12'h7A8;
        15'h1BCB: data = 12'h785;
        15'h1BCC: data = 12'h763;
        15'h1BCD: data = 12'h77B;
        15'h1BCE: data = 12'h798;
        15'h1BCF: data = 12'h7D0;
        15'h1BD0: data = 12'h338;
        15'h1BD1: data = 12'h0DC;
        15'h1BD2: data = 12'h151;
        15'h1BD3: data = 12'h1E2;
        15'h1BD4: data = 12'h281;
        15'h1BD5: data = 12'h33C;
        15'h1BD6: data = 12'h3F9;
        15'h1BD7: data = 12'h4C7;
        15'h1BD8: data = 12'h50D;
        15'h1BD9: data = 12'h682;
        15'h1BDA: data = 12'h773;
        15'h1BDB: data = 12'h0FD;
        15'h1BDC: data = 12'h1A3;
        15'h1BDD: data = 12'h2C7;
        15'h1BDE: data = 12'h3E1;
        15'h1BDF: data = 12'h505;
        15'h1BE0: data = 12'h61E;
        15'h1BE1: data = 12'h73A;
        15'h1BE2: data = 12'h559;
        15'h1BE3: data = 12'h1C1;
        15'h1BE4: data = 12'h2D7;
        15'h1BE5: data = 12'h3EF;
        15'h1BE6: data = 12'h502;
        15'h1BE7: data = 12'h60C;
        15'h1BE8: data = 12'h712;
        15'h1BE9: data = 12'h806;
        15'h1BEA: data = 12'h132;
        15'h1BEB: data = 12'h204;
        15'h1BEC: data = 12'h2CF;
        15'h1BED: data = 12'h384;
        15'h1BEE: data = 12'h429;
        15'h1BEF: data = 12'h4B4;
        15'h1BF0: data = 12'h542;
        15'h1BF1: data = 12'h5AA;
        15'h1BF2: data = 12'h5F9;
        15'h1BF3: data = 12'h64E;
        15'h1BF4: data = 12'h675;
        15'h1BF5: data = 12'h696;
        15'h1BF6: data = 12'h698;
        15'h1BF7: data = 12'h50D;
        15'h1BF8: data = 12'h657;
        15'h1BF9: data = 12'h613;
        15'h1BFA: data = 12'h5BC;
        15'h1BFB: data = 12'h54E;
        15'h1BFC: data = 12'h4CB;
        15'h1BFD: data = 12'h436;
        15'h1BFE: data = 12'h391;
        15'h1BFF: data = 12'h2E1;
        15'h1C00: data = 12'h21C;
        15'h1C01: data = 12'h14D;
        15'h1C02: data = 12'h071;
        15'h1C03: data = 12'h742;
        15'h1C04: data = 12'h641;
        15'h1C05: data = 12'h53C;
        15'h1C06: data = 12'h423;
        15'h1C07: data = 12'h312;
        15'h1C08: data = 12'h1EC;
        15'h1C09: data = 12'h0C9;
        15'h1C0A: data = 12'h763;
        15'h1C0B: data = 12'h63D;
        15'h1C0C: data = 12'h520;
        15'h1C0D: data = 12'h40F;
        15'h1C0E: data = 12'h2F5;
        15'h1C0F: data = 12'h1E1;
        15'h1C10: data = 12'h0DB;
        15'h1C11: data = 12'h7A9;
        15'h1C12: data = 12'h6AF;
        15'h1C13: data = 12'h5C2;
        15'h1C14: data = 12'h4E4;
        15'h1C15: data = 12'h40E;
        15'h1C16: data = 12'h50D;
        15'h1C17: data = 12'h28E;
        15'h1C18: data = 12'h1F2;
        15'h1C19: data = 12'h164;
        15'h1C1A: data = 12'h0FD;
        15'h1C1B: data = 12'h09D;
        15'h1C1C: data = 12'h04A;
        15'h1C1D: data = 12'h7A4;
        15'h1C1E: data = 12'h786;
        15'h1C1F: data = 12'h764;
        15'h1C20: data = 12'h782;
        15'h1C21: data = 12'h781;
        15'h1C22: data = 12'h7B4;
        15'h1C23: data = 12'h7F7;
        15'h1C24: data = 12'h0B2;
        15'h1C25: data = 12'h122;
        15'h1C26: data = 12'h1B0;
        15'h1C27: data = 12'h255;
        15'h1C28: data = 12'h2FF;
        15'h1C29: data = 12'h3B9;
        15'h1C2A: data = 12'h485;
        15'h1C2B: data = 12'h54D;
        15'h1C2C: data = 12'h636;
        15'h1C2D: data = 12'h71E;
        15'h1C2E: data = 12'h817;
        15'h1C2F: data = 12'h150;
        15'h1C30: data = 12'h260;
        15'h1C31: data = 12'h382;
        15'h1C32: data = 12'h4A4;
        15'h1C33: data = 12'h5BF;
        15'h1C34: data = 12'h6E9;
        15'h1C35: data = 12'h50D;
        15'h1C36: data = 12'h163;
        15'h1C37: data = 12'h285;
        15'h1C38: data = 12'h397;
        15'h1C39: data = 12'h4AD;
        15'h1C3A: data = 12'h5AA;
        15'h1C3B: data = 12'h6B9;
        15'h1C3C: data = 12'h7B1;
        15'h1C3D: data = 12'h0E1;
        15'h1C3E: data = 12'h1BE;
        15'h1C3F: data = 12'h290;
        15'h1C40: data = 12'h348;
        15'h1C41: data = 12'h3FC;
        15'h1C42: data = 12'h49A;
        15'h1C43: data = 12'h510;
        15'h1C44: data = 12'h581;
        15'h1C45: data = 12'h5E6;
        15'h1C46: data = 12'h627;
        15'h1C47: data = 12'h66D;
        15'h1C48: data = 12'h692;
        15'h1C49: data = 12'h698;
        15'h1C4A: data = 12'h696;
        15'h1C4B: data = 12'h66D;
        15'h1C4C: data = 12'h636;
        15'h1C4D: data = 12'h5D8;
        15'h1C4E: data = 12'h56C;
        15'h1C4F: data = 12'h4F7;
        15'h1C50: data = 12'h46C;
        15'h1C51: data = 12'h3D5;
        15'h1C52: data = 12'h322;
        15'h1C53: data = 12'h265;
        15'h1C54: data = 12'h50D;
        15'h1C55: data = 12'h0BD;
        15'h1C56: data = 12'h78E;
        15'h1C57: data = 12'h699;
        15'h1C58: data = 12'h592;
        15'h1C59: data = 12'h48B;
        15'h1C5A: data = 12'h368;
        15'h1C5B: data = 12'h24C;
        15'h1C5C: data = 12'h12D;
        15'h1C5D: data = 12'h02A;
        15'h1C5E: data = 12'h6A0;
        15'h1C5F: data = 12'h57B;
        15'h1C60: data = 12'h468;
        15'h1C61: data = 12'h34F;
        15'h1C62: data = 12'h23D;
        15'h1C63: data = 12'h12C;
        15'h1C64: data = 12'h031;
        15'h1C65: data = 12'h701;
        15'h1C66: data = 12'h60F;
        15'h1C67: data = 12'h52A;
        15'h1C68: data = 12'h457;
        15'h1C69: data = 12'h38A;
        15'h1C6A: data = 12'h2CF;
        15'h1C6B: data = 12'h227;
        15'h1C6C: data = 12'h191;
        15'h1C6D: data = 12'h10C;
        15'h1C6E: data = 12'h0BE;
        15'h1C6F: data = 12'h063;
        15'h1C70: data = 12'h6EA;
        15'h1C71: data = 12'h786;
        15'h1C72: data = 12'h774;
        15'h1C73: data = 12'h50D;
        15'h1C74: data = 12'h77B;
        15'h1C75: data = 12'h79E;
        15'h1C76: data = 12'h7E7;
        15'h1C77: data = 12'h096;
        15'h1C78: data = 12'h101;
        15'h1C79: data = 12'h179;
        15'h1C7A: data = 12'h210;
        15'h1C7B: data = 12'h2B9;
        15'h1C7C: data = 12'h377;
        15'h1C7D: data = 12'h43C;
        15'h1C7E: data = 12'h50B;
        15'h1C7F: data = 12'h5EB;
        15'h1C80: data = 12'h6DC;
        15'h1C81: data = 12'h7CC;
        15'h1C82: data = 12'h0FF;
        15'h1C83: data = 12'h205;
        15'h1C84: data = 12'h316;
        15'h1C85: data = 12'h43C;
        15'h1C86: data = 12'h557;
        15'h1C87: data = 12'h684;
        15'h1C88: data = 12'h7A5;
        15'h1C89: data = 12'h10D;
        15'h1C8A: data = 12'h226;
        15'h1C8B: data = 12'h33B;
        15'h1C8C: data = 12'h44D;
        15'h1C8D: data = 12'h557;
        15'h1C8E: data = 12'h660;
        15'h1C8F: data = 12'h75D;
        15'h1C90: data = 12'h177;
        15'h1C91: data = 12'h177;
        15'h1C92: data = 12'h50D;
        15'h1C93: data = 12'h30E;
        15'h1C94: data = 12'h3C0;
        15'h1C95: data = 12'h461;
        15'h1C96: data = 12'h4EF;
        15'h1C97: data = 12'h55A;
        15'h1C98: data = 12'h5C6;
        15'h1C99: data = 12'h608;
        15'h1C9A: data = 12'h64A;
        15'h1C9B: data = 12'h689;
        15'h1C9C: data = 12'h694;
        15'h1C9D: data = 12'h698;
        15'h1C9E: data = 12'h679;
        15'h1C9F: data = 12'h63D;
        15'h1CA0: data = 12'h5F1;
        15'h1CA1: data = 12'h592;
        15'h1CA2: data = 12'h52A;
        15'h1CA3: data = 12'h498;
        15'h1CA4: data = 12'h400;
        15'h1CA5: data = 12'h355;
        15'h1CA6: data = 12'h29E;
        15'h1CA7: data = 12'h1D5;
        15'h1CA8: data = 12'h105;
        15'h1CA9: data = 12'h255;
        15'h1CAA: data = 12'h6ED;
        15'h1CAB: data = 12'h5EE;
        15'h1CAC: data = 12'h4E4;
        15'h1CAD: data = 12'h3CC;
        15'h1CAE: data = 12'h2AA;
        15'h1CAF: data = 12'h18B;
        15'h1CB0: data = 12'h06B;
        15'h1CB1: data = 12'h50D;
        15'h1CB2: data = 12'h5D9;
        15'h1CB3: data = 12'h4C5;
        15'h1CB4: data = 12'h3A5;
        15'h1CB5: data = 12'h299;
        15'h1CB6: data = 12'h189;
        15'h1CB7: data = 12'h086;
        15'h1CB8: data = 12'h74F;
        15'h1CB9: data = 12'h665;
        15'h1CBA: data = 12'h574;
        15'h1CBB: data = 12'h49B;
        15'h1CBC: data = 12'h3C7;
        15'h1CBD: data = 12'h307;
        15'h1CBE: data = 12'h25C;
        15'h1CBF: data = 12'h1C7;
        15'h1CC0: data = 12'h133;
        15'h1CC1: data = 12'h0D8;
        15'h1CC2: data = 12'h087;
        15'h1CC3: data = 12'h032;
        15'h1CC4: data = 12'h7AA;
        15'h1CC5: data = 12'h785;
        15'h1CC6: data = 12'h761;
        15'h1CC7: data = 12'h77D;
        15'h1CC8: data = 12'h796;
        15'h1CC9: data = 12'h7D2;
        15'h1CCA: data = 12'h39C;
        15'h1CCB: data = 12'h0DA;
        15'h1CCC: data = 12'h14A;
        15'h1CCD: data = 12'h1D8;
        15'h1CCE: data = 12'h276;
        15'h1CCF: data = 12'h334;
        15'h1CD0: data = 12'h50D;
        15'h1CD1: data = 12'h4C7;
        15'h1CD2: data = 12'h5A1;
        15'h1CD3: data = 12'h688;
        15'h1CD4: data = 12'h772;
        15'h1CD5: data = 12'h11C;
        15'h1CD6: data = 12'h1A1;
        15'h1CD7: data = 12'h2C0;
        15'h1CD8: data = 12'h3D9;
        15'h1CD9: data = 12'h4FF;
        15'h1CDA: data = 12'h61F;
        15'h1CDB: data = 12'h736;
        15'h1CDC: data = 12'h57A;
        15'h1CDD: data = 12'h1C5;
        15'h1CDE: data = 12'h2DE;
        15'h1CDF: data = 12'h3F5;
        15'h1CE0: data = 12'h500;
        15'h1CE1: data = 12'h60C;
        15'h1CE2: data = 12'h70E;
        15'h1CE3: data = 12'h7FF;
        15'h1CE4: data = 12'h12C;
        15'h1CE5: data = 12'h1FD;
        15'h1CE6: data = 12'h2D2;
        15'h1CE7: data = 12'h385;
        15'h1CE8: data = 12'h42A;
        15'h1CE9: data = 12'h4B7;
        15'h1CEA: data = 12'h53B;
        15'h1CEB: data = 12'h5A3;
        15'h1CEC: data = 12'h5F4;
        15'h1CED: data = 12'h648;
        15'h1CEE: data = 12'h66B;
        15'h1CEF: data = 12'h50D;
        15'h1CF0: data = 12'h694;
        15'h1CF1: data = 12'h677;
        15'h1CF2: data = 12'h654;
        15'h1CF3: data = 12'h60E;
        15'h1CF4: data = 12'h5B5;
        15'h1CF5: data = 12'h54C;
        15'h1CF6: data = 12'h4CA;
        15'h1CF7: data = 12'h438;
        15'h1CF8: data = 12'h390;
        15'h1CF9: data = 12'h2DC;
        15'h1CFA: data = 12'h219;
        15'h1CFB: data = 12'h146;
        15'h1CFC: data = 12'h06B;
        15'h1CFD: data = 12'h73D;
        15'h1CFE: data = 12'h63F;
        15'h1CFF: data = 12'h53A;
        15'h1D00: data = 12'h426;
        15'h1D01: data = 12'h310;
        15'h1D02: data = 12'h1EE;
        15'h1D03: data = 12'h0CA;
        15'h1D04: data = 12'h760;
        15'h1D05: data = 12'h639;
        15'h1D06: data = 12'h51B;
        15'h1D07: data = 12'h406;
        15'h1D08: data = 12'h2F0;
        15'h1D09: data = 12'h1DC;
        15'h1D0A: data = 12'h0D8;
        15'h1D0B: data = 12'h775;
        15'h1D0C: data = 12'h6AE;
        15'h1D0D: data = 12'h5C2;
        15'h1D0E: data = 12'h50D;
        15'h1D0F: data = 12'h40C;
        15'h1D10: data = 12'h344;
        15'h1D11: data = 12'h28D;
        15'h1D12: data = 12'h1F1;
        15'h1D13: data = 12'h166;
        15'h1D14: data = 12'h0FD;
        15'h1D15: data = 12'h09A;
        15'h1D16: data = 12'h045;
        15'h1D17: data = 12'h7A5;
        15'h1D18: data = 12'h787;
        15'h1D19: data = 12'h766;
        15'h1D1A: data = 12'h77E;
        15'h1D1B: data = 12'h783;
        15'h1D1C: data = 12'h7B4;
        15'h1D1D: data = 12'h7F2;
        15'h1D1E: data = 12'h0B4;
        15'h1D1F: data = 12'h11C;
        15'h1D20: data = 12'h1AE;
        15'h1D21: data = 12'h24E;
        15'h1D22: data = 12'h2F9;
        15'h1D23: data = 12'h3B5;
        15'h1D24: data = 12'h488;
        15'h1D25: data = 12'h551;
        15'h1D26: data = 12'h63C;
        15'h1D27: data = 12'h724;
        15'h1D28: data = 12'h81C;
        15'h1D29: data = 12'h151;
        15'h1D2A: data = 12'h25E;
        15'h1D2B: data = 12'h376;
        15'h1D2C: data = 12'h49C;
        15'h1D2D: data = 12'h50D;
        15'h1D2E: data = 12'h6EB;
        15'h1D2F: data = 12'h801;
        15'h1D30: data = 12'h167;
        15'h1D31: data = 12'h289;
        15'h1D32: data = 12'h398;
        15'h1D33: data = 12'h4AD;
        15'h1D34: data = 12'h5AE;
        15'h1D35: data = 12'h6B9;
        15'h1D36: data = 12'h7AE;
        15'h1D37: data = 12'h0DF;
        15'h1D38: data = 12'h1C2;
        15'h1D39: data = 12'h291;
        15'h1D3A: data = 12'h346;
        15'h1D3B: data = 12'h3F7;
        15'h1D3C: data = 12'h495;
        15'h1D3D: data = 12'h518;
        15'h1D3E: data = 12'h587;
        15'h1D3F: data = 12'h5EA;
        15'h1D40: data = 12'h62A;
        15'h1D41: data = 12'h667;
        15'h1D42: data = 12'h686;
        15'h1D43: data = 12'h68F;
        15'h1D44: data = 12'h693;
        15'h1D45: data = 12'h66A;
        15'h1D46: data = 12'h635;
        15'h1D47: data = 12'h5D7;
        15'h1D48: data = 12'h572;
        15'h1D49: data = 12'h4FE;
        15'h1D4A: data = 12'h46F;
        15'h1D4B: data = 12'h3CB;
        15'h1D4C: data = 12'h50D;
        15'h1D4D: data = 12'h25C;
        15'h1D4E: data = 12'h18E;
        15'h1D4F: data = 12'h0B4;
        15'h1D50: data = 12'h78E;
        15'h1D51: data = 12'h698;
        15'h1D52: data = 12'h596;
        15'h1D53: data = 12'h48B;
        15'h1D54: data = 12'h370;
        15'h1D55: data = 12'h254;
        15'h1D56: data = 12'h12F;
        15'h1D57: data = 12'h01A;
        15'h1D58: data = 12'h69F;
        15'h1D59: data = 12'h579;
        15'h1D5A: data = 12'h464;
        15'h1D5B: data = 12'h345;
        15'h1D5C: data = 12'h236;
        15'h1D5D: data = 12'h127;
        15'h1D5E: data = 12'h0A5;
        15'h1D5F: data = 12'h6FE;
        15'h1D60: data = 12'h611;
        15'h1D61: data = 12'h530;
        15'h1D62: data = 12'h460;
        15'h1D63: data = 12'h38D;
        15'h1D64: data = 12'h2D4;
        15'h1D65: data = 12'h227;
        15'h1D66: data = 12'h18F;
        15'h1D67: data = 12'h10B;
        15'h1D68: data = 12'h0B1;
        15'h1D69: data = 12'h060;
        15'h1D6A: data = 12'h7C5;
        15'h1D6B: data = 12'h50D;
        15'h1D6C: data = 12'h776;
        15'h1D6D: data = 12'h761;
        15'h1D6E: data = 12'h782;
        15'h1D6F: data = 12'h7A8;
        15'h1D70: data = 12'h7E8;
        15'h1D71: data = 12'h095;
        15'h1D72: data = 12'h0FF;
        15'h1D73: data = 12'h175;
        15'h1D74: data = 12'h206;
        15'h1D75: data = 12'h2B0;
        15'h1D76: data = 12'h36B;
        15'h1D77: data = 12'h43A;
        15'h1D78: data = 12'h50F;
        15'h1D79: data = 12'h5F6;
        15'h1D7A: data = 12'h6E5;
        15'h1D7B: data = 12'h7D5;
        15'h1D7C: data = 12'h102;
        15'h1D7D: data = 12'h204;
        15'h1D7E: data = 12'h30D;
        15'h1D7F: data = 12'h432;
        15'h1D80: data = 12'h54E;
        15'h1D81: data = 12'h67A;
        15'h1D82: data = 12'h7A2;
        15'h1D83: data = 12'h111;
        15'h1D84: data = 12'h225;
        15'h1D85: data = 12'h343;
        15'h1D86: data = 12'h45A;
        15'h1D87: data = 12'h560;
        15'h1D88: data = 12'h664;
        15'h1D89: data = 12'h75F;
        15'h1D8A: data = 12'h50D;
        15'h1D8B: data = 12'h16F;
        15'h1D8C: data = 12'h245;
        15'h1D8D: data = 12'h30F;
        15'h1D8E: data = 12'h3C1;
        15'h1D8F: data = 12'h464;
        15'h1D90: data = 12'h4F9;
        15'h1D91: data = 12'h56B;
        15'h1D92: data = 12'h5D0;
        15'h1D93: data = 12'h605;
        15'h1D94: data = 12'h643;
        15'h1D95: data = 12'h67D;
        15'h1D96: data = 12'h681;
        15'h1D97: data = 12'h689;
        15'h1D98: data = 12'h671;
        15'h1D99: data = 12'h63F;
        15'h1D9A: data = 12'h5F4;
        15'h1D9B: data = 12'h59C;
        15'h1D9C: data = 12'h534;
        15'h1D9D: data = 12'h4A1;
        15'h1D9E: data = 12'h407;
        15'h1D9F: data = 12'h358;
        15'h1DA0: data = 12'h29D;
        15'h1DA1: data = 12'h1CC;
        15'h1DA2: data = 12'h0F4;
        15'h1DA3: data = 12'h109;
        15'h1DA4: data = 12'h6E6;
        15'h1DA5: data = 12'h5EC;
        15'h1DA6: data = 12'h4E0;
        15'h1DA7: data = 12'h3CD;
        15'h1DA8: data = 12'h2B2;
        15'h1DA9: data = 12'h50D;
        15'h1DAA: data = 12'h078;
        15'h1DAB: data = 12'h6FC;
        15'h1DAC: data = 12'h5DF;
        15'h1DAD: data = 12'h4C5;
        15'h1DAE: data = 12'h39F;
        15'h1DAF: data = 12'h28A;
        15'h1DB0: data = 12'h178;
        15'h1DB1: data = 12'h076;
        15'h1DB2: data = 12'h745;
        15'h1DB3: data = 12'h660;
        15'h1DB4: data = 12'h576;
        15'h1DB5: data = 12'h49F;
        15'h1DB6: data = 12'h3D9;
        15'h1DB7: data = 12'h31D;
        15'h1DB8: data = 12'h26B;
        15'h1DB9: data = 12'h1CE;
        15'h1DBA: data = 12'h131;
        15'h1DBB: data = 12'h0D2;
        15'h1DBC: data = 12'h077;
        15'h1DBD: data = 12'h02B;
        15'h1DBE: data = 12'h79C;
        15'h1DBF: data = 12'h780;
        15'h1DC0: data = 12'h764;
        15'h1DC1: data = 12'h785;
        15'h1DC2: data = 12'h7A4;
        15'h1DC3: data = 12'h7E0;
        15'h1DC4: data = 12'h731;
        15'h1DC5: data = 12'h0DD;
        15'h1DC6: data = 12'h14B;
        15'h1DC7: data = 12'h1CE;
        15'h1DC8: data = 12'h50D;
        15'h1DC9: data = 12'h329;
        15'h1DCA: data = 12'h3E9;
        15'h1DCB: data = 12'h4C1;
        15'h1DCC: data = 12'h59C;
        15'h1DCD: data = 12'h68F;
        15'h1DCE: data = 12'h783;
        15'h1DCF: data = 12'h0A9;
        15'h1DD0: data = 12'h1B4;
        15'h1DD1: data = 12'h2C6;
        15'h1DD2: data = 12'h3D6;
        15'h1DD3: data = 12'h4F3;
        15'h1DD4: data = 12'h610;
        15'h1DD5: data = 12'h729;
        15'h1DD6: data = 12'h2BC;
        15'h1DD7: data = 12'h1C3;
        15'h1DD8: data = 12'h2E7;
        15'h1DD9: data = 12'h403;
        15'h1DDA: data = 12'h516;
        15'h1DDB: data = 12'h617;
        15'h1DDC: data = 12'h70C;
        15'h1DDD: data = 12'h7FA;
        15'h1DDE: data = 12'h11A;
        15'h1DDF: data = 12'h1F3;
        15'h1DE0: data = 12'h2BD;
        15'h1DE1: data = 12'h380;
        15'h1DE2: data = 12'h42F;
        15'h1DE3: data = 12'h4C1;
        15'h1DE4: data = 12'h549;
        15'h1DE5: data = 12'h5B7;
        15'h1DE6: data = 12'h603;
        15'h1DE7: data = 12'h50D;
        15'h1DE8: data = 12'h66D;
        15'h1DE9: data = 12'h686;
        15'h1DEA: data = 12'h686;
        15'h1DEB: data = 12'h665;
        15'h1DEC: data = 12'h649;
        15'h1DED: data = 12'h610;
        15'h1DEE: data = 12'h5BF;
        15'h1DEF: data = 12'h560;
        15'h1DF0: data = 12'h4E2;
        15'h1DF1: data = 12'h44B;
        15'h1DF2: data = 12'h39C;
        15'h1DF3: data = 12'h2E5;
        15'h1DF4: data = 12'h217;
        15'h1DF5: data = 12'h13E;
        15'h1DF6: data = 12'h05E;
        15'h1DF7: data = 12'h72F;
        15'h1DF8: data = 12'h633;
        15'h1DF9: data = 12'h532;
        15'h1DFA: data = 12'h423;
        15'h1DFB: data = 12'h317;
        15'h1DFC: data = 12'h1F9;
        15'h1DFD: data = 12'h0D9;
        15'h1DFE: data = 12'h76A;
        15'h1DFF: data = 12'h64E;
        15'h1E00: data = 12'h526;
        15'h1E01: data = 12'h40C;
        15'h1E02: data = 12'h2ED;
        15'h1E03: data = 12'h1D1;
        15'h1E04: data = 12'h0C9;
        15'h1E05: data = 12'h7A2;
        15'h1E06: data = 12'h50D;
        15'h1E07: data = 12'h5BD;
        15'h1E08: data = 12'h4EB;
        15'h1E09: data = 12'h416;
        15'h1E0A: data = 12'h355;
        15'h1E0B: data = 12'h2A0;
        15'h1E0C: data = 12'h200;
        15'h1E0D: data = 12'h171;
        15'h1E0E: data = 12'h0FB;
        15'h1E0F: data = 12'h092;
        15'h1E10: data = 12'h038;
        15'h1E11: data = 12'h793;
        15'h1E12: data = 12'h774;
        15'h1E13: data = 12'h75A;
        15'h1E14: data = 12'h77F;
        15'h1E15: data = 12'h787;
        15'h1E16: data = 12'h7C5;
        15'h1E17: data = 12'h809;
        15'h1E18: data = 12'h0C4;
        15'h1E19: data = 12'h12D;
        15'h1E1A: data = 12'h1AF;
        15'h1E1B: data = 12'h242;
        15'h1E1C: data = 12'h2EB;
        15'h1E1D: data = 12'h3A4;
        15'h1E1E: data = 12'h476;
        15'h1E1F: data = 12'h549;
        15'h1E20: data = 12'h63C;
        15'h1E21: data = 12'h72C;
        15'h1E22: data = 12'h82E;
        15'h1E23: data = 12'h160;
        15'h1E24: data = 12'h272;
        15'h1E25: data = 12'h50D;
        15'h1E26: data = 12'h49B;
        15'h1E27: data = 12'h5B1;
        15'h1E28: data = 12'h6D5;
        15'h1E29: data = 12'h7ED;
        15'h1E2A: data = 12'h157;
        15'h1E2B: data = 12'h285;
        15'h1E2C: data = 12'h39B;
        15'h1E2D: data = 12'h4BA;
        15'h1E2E: data = 12'h5C0;
        15'h1E2F: data = 12'h6CD;
        15'h1E30: data = 12'h7B7;
        15'h1E31: data = 12'h0DF;
        15'h1E32: data = 12'h1B4;
        15'h1E33: data = 12'h282;
        15'h1E34: data = 12'h339;
        15'h1E35: data = 12'h3F0;
        15'h1E36: data = 12'h494;
        15'h1E37: data = 12'h51C;
        15'h1E38: data = 12'h593;
        15'h1E39: data = 12'h5FA;
        15'h1E3A: data = 12'h639;
        15'h1E3B: data = 12'h679;
        15'h1E3C: data = 12'h694;
        15'h1E3D: data = 12'h68D;
        15'h1E3E: data = 12'h688;
        15'h1E3F: data = 12'h65F;
        15'h1E40: data = 12'h628;
        15'h1E41: data = 12'h5CC;
        15'h1E42: data = 12'h56D;
        15'h1E43: data = 12'h507;
        15'h1E44: data = 12'h50D;
        15'h1E45: data = 12'h3E2;
        15'h1E46: data = 12'h330;
        15'h1E47: data = 12'h269;
        15'h1E48: data = 12'h196;
        15'h1E49: data = 12'h0B3;
        15'h1E4A: data = 12'h782;
        15'h1E4B: data = 12'h688;
        15'h1E4C: data = 12'h580;
        15'h1E4D: data = 12'h47A;
        15'h1E4E: data = 12'h361;
        15'h1E4F: data = 12'h24B;
        15'h1E50: data = 12'h13A;
        15'h1E51: data = 12'h1EC;
        15'h1E52: data = 12'h6AE;
        15'h1E53: data = 12'h58B;
        15'h1E54: data = 12'h473;
        15'h1E55: data = 12'h352;
        15'h1E56: data = 12'h239;
        15'h1E57: data = 12'h11F;
        15'h1E58: data = 12'h020;
        15'h1E59: data = 12'h6F1;
        15'h1E5A: data = 12'h602;
        15'h1E5B: data = 12'h523;
        15'h1E5C: data = 12'h458;
        15'h1E5D: data = 12'h38E;
        15'h1E5E: data = 12'h2DE;
        15'h1E5F: data = 12'h23A;
        15'h1E60: data = 12'h1A2;
        15'h1E61: data = 12'h121;
        15'h1E62: data = 12'h0C1;
        15'h1E63: data = 12'h50D;
        15'h1E64: data = 12'h7AE;
        15'h1E65: data = 12'h771;
        15'h1E66: data = 12'h75F;
        15'h1E67: data = 12'h755;
        15'h1E68: data = 12'h775;
        15'h1E69: data = 12'h7A7;
        15'h1E6A: data = 12'h7F6;
        15'h1E6B: data = 12'h0B6;
        15'h1E6C: data = 12'h113;
        15'h1E6D: data = 12'h182;
        15'h1E6E: data = 12'h217;
        15'h1E6F: data = 12'h2B4;
        15'h1E70: data = 12'h368;
        15'h1E71: data = 12'h42A;
        15'h1E72: data = 12'h4FD;
        15'h1E73: data = 12'h5E2;
        15'h1E74: data = 12'h6DA;
        15'h1E75: data = 12'h7D4;
        15'h1E76: data = 12'h10C;
        15'h1E77: data = 12'h216;
        15'h1E78: data = 12'h324;
        15'h1E79: data = 12'h445;
        15'h1E7A: data = 12'h55B;
        15'h1E7B: data = 12'h67B;
        15'h1E7C: data = 12'h795;
        15'h1E7D: data = 12'h100;
        15'h1E7E: data = 12'h216;
        15'h1E7F: data = 12'h339;
        15'h1E80: data = 12'h458;
        15'h1E81: data = 12'h56B;
        15'h1E82: data = 12'h50D;
        15'h1E83: data = 12'h76C;
        15'h1E84: data = 12'h3F3;
        15'h1E85: data = 12'h175;
        15'h1E86: data = 12'h248;
        15'h1E87: data = 12'h304;
        15'h1E88: data = 12'h3B3;
        15'h1E89: data = 12'h452;
        15'h1E8A: data = 12'h4E9;
        15'h1E8B: data = 12'h563;
        15'h1E8C: data = 12'h5D3;
        15'h1E8D: data = 12'h618;
        15'h1E8E: data = 12'h654;
        15'h1E8F: data = 12'h68E;
        15'h1E90: data = 12'h691;
        15'h1E91: data = 12'h692;
        15'h1E92: data = 12'h667;
        15'h1E93: data = 12'h62F;
        15'h1E94: data = 12'h5E2;
        15'h1E95: data = 12'h588;
        15'h1E96: data = 12'h52A;
        15'h1E97: data = 12'h49D;
        15'h1E98: data = 12'h409;
        15'h1E99: data = 12'h363;
        15'h1E9A: data = 12'h2AB;
        15'h1E9B: data = 12'h1E5;
        15'h1E9C: data = 12'h105;
        15'h1E9D: data = 12'h021;
        15'h1E9E: data = 12'h6E3;
        15'h1E9F: data = 12'h5DB;
        15'h1EA0: data = 12'h4CB;
        15'h1EA1: data = 12'h50D;
        15'h1EA2: data = 12'h2A1;
        15'h1EA3: data = 12'h18A;
        15'h1EA4: data = 12'h073;
        15'h1EA5: data = 12'h702;
        15'h1EA6: data = 12'h5EC;
        15'h1EA7: data = 12'h4D4;
        15'h1EA8: data = 12'h3AC;
        15'h1EA9: data = 12'h29C;
        15'h1EAA: data = 12'h185;
        15'h1EAB: data = 12'h07E;
        15'h1EAC: data = 12'h744;
        15'h1EAD: data = 12'h657;
        15'h1EAE: data = 12'h565;
        15'h1EAF: data = 12'h491;
        15'h1EB0: data = 12'h3C4;
        15'h1EB1: data = 12'h30E;
        15'h1EB2: data = 12'h265;
        15'h1EB3: data = 12'h1D6;
        15'h1EB4: data = 12'h147;
        15'h1EB5: data = 12'h0E7;
        15'h1EB6: data = 12'h084;
        15'h1EB7: data = 12'h02E;
        15'h1EB8: data = 12'h79F;
        15'h1EB9: data = 12'h77D;
        15'h1EBA: data = 12'h755;
        15'h1EBB: data = 12'h770;
        15'h1EBC: data = 12'h792;
        15'h1EBD: data = 12'h7D2;
        15'h1EBE: data = 12'h296;
        15'h1EBF: data = 12'h0E3;
        15'h1EC0: data = 12'h50D;
        15'h1EC1: data = 12'h1E5;
        15'h1EC2: data = 12'h284;
        15'h1EC3: data = 12'h337;
        15'h1EC4: data = 12'h3EE;
        15'h1EC5: data = 12'h4BD;
        15'h1EC6: data = 12'h590;
        15'h1EC7: data = 12'h67E;
        15'h1EC8: data = 12'h76E;
        15'h1EC9: data = 12'h0DF;
        15'h1ECA: data = 12'h1AB;
        15'h1ECB: data = 12'h2D0;
        15'h1ECC: data = 12'h3E7;
        15'h1ECD: data = 12'h508;
        15'h1ECE: data = 12'h625;
        15'h1ECF: data = 12'h73A;
        15'h1ED0: data = 12'h40B;
        15'h1ED1: data = 12'h1BC;
        15'h1ED2: data = 12'h2D5;
        15'h1ED3: data = 12'h3F2;
        15'h1ED4: data = 12'h506;
        15'h1ED5: data = 12'h617;
        15'h1ED6: data = 12'h71B;
        15'h1ED7: data = 12'h80D;
        15'h1ED8: data = 12'h12D;
        15'h1ED9: data = 12'h204;
        15'h1EDA: data = 12'h2C9;
        15'h1EDB: data = 12'h37B;
        15'h1EDC: data = 12'h424;
        15'h1EDD: data = 12'h4B3;
        15'h1EDE: data = 12'h53D;
        15'h1EDF: data = 12'h50D;
        15'h1EE0: data = 12'h5FA;
        15'h1EE1: data = 12'h654;
        15'h1EE2: data = 12'h677;
        15'h1EE3: data = 12'h697;
        15'h1EE4: data = 12'h695;
        15'h1EE5: data = 12'h671;
        15'h1EE6: data = 12'h655;
        15'h1EE7: data = 12'h60D;
        15'h1EE8: data = 12'h5AD;
        15'h1EE9: data = 12'h54A;
        15'h1EEA: data = 12'h4CD;
        15'h1EEB: data = 12'h43A;
        15'h1EEC: data = 12'h390;
        15'h1EED: data = 12'h2E3;
        15'h1EEE: data = 12'h221;
        15'h1EEF: data = 12'h151;
        15'h1EF0: data = 12'h06D;
        15'h1EF1: data = 12'h73B;
        15'h1EF2: data = 12'h63C;
        15'h1EF3: data = 12'h538;
        15'h1EF4: data = 12'h41E;
        15'h1EF5: data = 12'h30C;
        15'h1EF6: data = 12'h1E8;
        15'h1EF7: data = 12'h0C9;
        15'h1EF8: data = 12'h762;
        15'h1EF9: data = 12'h63E;
        15'h1EFA: data = 12'h51F;
        15'h1EFB: data = 12'h414;
        15'h1EFC: data = 12'h2F8;
        15'h1EFD: data = 12'h1E3;
        15'h1EFE: data = 12'h50D;
        15'h1EFF: data = 12'h7A0;
        15'h1F00: data = 12'h6AC;
        15'h1F01: data = 12'h5BC;
        15'h1F02: data = 12'h4DE;
        15'h1F03: data = 12'h40B;
        15'h1F04: data = 12'h346;
        15'h1F05: data = 12'h291;
        15'h1F06: data = 12'h1F3;
        15'h1F07: data = 12'h16E;
        15'h1F08: data = 12'h102;
        15'h1F09: data = 12'h09C;
        15'h1F0A: data = 12'h047;
        15'h1F0B: data = 12'h7A1;
        15'h1F0C: data = 12'h782;
        15'h1F0D: data = 12'h762;
        15'h1F0E: data = 12'h77F;
        15'h1F0F: data = 12'h780;
        15'h1F10: data = 12'h7AF;
        15'h1F11: data = 12'h7F3;
        15'h1F12: data = 12'h0B6;
        15'h1F13: data = 12'h128;
        15'h1F14: data = 12'h1B4;
        15'h1F15: data = 12'h257;
        15'h1F16: data = 12'h2FB;
        15'h1F17: data = 12'h3B7;
        15'h1F18: data = 12'h486;
        15'h1F19: data = 12'h54C;
        15'h1F1A: data = 12'h637;
        15'h1F1B: data = 12'h723;
        15'h1F1C: data = 12'h81C;
        15'h1F1D: data = 12'h50D;
        15'h1F1E: data = 12'h265;
        15'h1F1F: data = 12'h383;
        15'h1F20: data = 12'h4A4;
        15'h1F21: data = 12'h5B8;
        15'h1F22: data = 12'h6E4;
        15'h1F23: data = 12'h800;
        15'h1F24: data = 12'h165;
        15'h1F25: data = 12'h27D;
        15'h1F26: data = 12'h398;
        15'h1F27: data = 12'h4A9;
        15'h1F28: data = 12'h5AF;
        15'h1F29: data = 12'h6C1;
        15'h1F2A: data = 12'h7B5;
        15'h1F2B: data = 12'h0E9;
        15'h1F2C: data = 12'h1C1;
        15'h1F2D: data = 12'h292;
        15'h1F2E: data = 12'h347;
        15'h1F2F: data = 12'h3F6;
        15'h1F30: data = 12'h490;
        15'h1F31: data = 12'h50F;
        15'h1F32: data = 12'h584;
        15'h1F33: data = 12'h5E9;
        15'h1F34: data = 12'h62C;
        15'h1F35: data = 12'h66F;
        15'h1F36: data = 12'h695;
        15'h1F37: data = 12'h695;
        15'h1F38: data = 12'h697;
        15'h1F39: data = 12'h66B;
        15'h1F3A: data = 12'h635;
        15'h1F3B: data = 12'h5D4;
        15'h1F3C: data = 12'h50D;
        15'h1F3D: data = 12'h4F4;
        15'h1F3E: data = 12'h46B;
        15'h1F3F: data = 12'h3CF;
        default: data = 12'h000;
    endcase
end

endmodule

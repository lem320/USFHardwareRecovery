module rom_good1 (
    input [14:0] address,
    output reg [11:0] data
);

always @(*) begin
    case (address)
        15'h0000: data = 12'h058;
        15'h0001: data = 12'h056;
        15'h0002: data = 12'h059;
        15'h0003: data = 12'h05A;
        15'h0004: data = 12'h060;
        15'h0005: data = 12'h064;
        15'h0006: data = 12'h065;
        15'h0007: data = 12'h064;
        15'h0008: data = 12'h062;
        15'h0009: data = 12'h064;
        15'h000A: data = 12'h05B;
        15'h000B: data = 12'h058;
        15'h000C: data = 12'h05B;
        15'h000D: data = 12'h05C;
        15'h000E: data = 12'h059;
        15'h000F: data = 12'h05D;
        15'h0010: data = 12'h062;
        15'h0011: data = 12'h064;
        15'h0012: data = 12'h067;
        15'h0013: data = 12'h064;
        15'h0014: data = 12'h063;
        15'h0015: data = 12'h060;
        15'h0016: data = 12'h05C;
        15'h0017: data = 12'h057;
        15'h0018: data = 12'h057;
        15'h0019: data = 12'h05C;
        15'h001A: data = 12'h05C;
        15'h001B: data = 12'h05C;
        15'h001C: data = 12'h062;
        15'h001D: data = 12'h068;
        15'h001E: data = 12'h068;
        15'h001F: data = 12'h062;
        15'h0020: data = 12'h05F;
        15'h0021: data = 12'h05D;
        15'h0022: data = 12'h057;
        15'h0023: data = 12'h05B;
        15'h0024: data = 12'h05A;
        15'h0025: data = 12'h059;
        15'h0026: data = 12'h05F;
        15'h0027: data = 12'h060;
        15'h0028: data = 12'h062;
        15'h0029: data = 12'h066;
        15'h002A: data = 12'h066;
        15'h002B: data = 12'h061;
        15'h002C: data = 12'h05C;
        15'h002D: data = 12'h05B;
        15'h002E: data = 12'h05D;
        15'h002F: data = 12'h05C;
        15'h0030: data = 12'h060;
        15'h0031: data = 12'h061;
        15'h0032: data = 12'h062;
        15'h0033: data = 12'h068;
        15'h0034: data = 12'h066;
        15'h0035: data = 12'h069;
        15'h0036: data = 12'h065;
        15'h0037: data = 12'h061;
        15'h0038: data = 12'h05A;
        15'h0039: data = 12'h059;
        15'h003A: data = 12'h059;
        15'h003B: data = 12'h038;
        15'h003C: data = 12'h03B;
        15'h003D: data = 12'h03F;
        15'h003E: data = 12'h041;
        15'h003F: data = 12'h047;
        15'h0040: data = 12'h043;
        15'h0041: data = 12'h044;
        15'h0042: data = 12'h040;
        15'h0043: data = 12'h03C;
        15'h0044: data = 12'h039;
        15'h0045: data = 12'h03A;
        15'h0046: data = 12'h036;
        15'h0047: data = 12'h03B;
        15'h0048: data = 12'h03F;
        15'h0049: data = 12'h041;
        15'h004A: data = 12'h045;
        15'h004B: data = 12'h043;
        15'h004C: data = 12'h044;
        15'h004D: data = 12'h040;
        15'h004E: data = 12'h03D;
        15'h004F: data = 12'h039;
        15'h0050: data = 12'h038;
        15'h0051: data = 12'h037;
        15'h0052: data = 12'h03A;
        15'h0053: data = 12'h03E;
        15'h0054: data = 12'h041;
        15'h0055: data = 12'h048;
        15'h0056: data = 12'h046;
        15'h0057: data = 12'h04A;
        15'h0058: data = 12'h047;
        15'h0059: data = 12'h045;
        15'h005A: data = 12'h03C;
        15'h005B: data = 12'h039;
        15'h005C: data = 12'h035;
        15'h005D: data = 12'h035;
        15'h005E: data = 12'h03F;
        15'h005F: data = 12'h042;
        15'h0060: data = 12'h047;
        15'h0061: data = 12'h048;
        15'h0062: data = 12'h044;
        15'h0063: data = 12'h046;
        15'h0064: data = 12'h040;
        15'h0065: data = 12'h03B;
        15'h0066: data = 12'h03A;
        15'h0067: data = 12'h037;
        15'h0068: data = 12'h03C;
        15'h0069: data = 12'h03A;
        15'h006A: data = 12'h03F;
        15'h006B: data = 12'h045;
        15'h006C: data = 12'h046;
        15'h006D: data = 12'h044;
        15'h006E: data = 12'h045;
        15'h006F: data = 12'h03F;
        15'h0070: data = 12'h036;
        15'h0071: data = 12'h806;
        15'h0072: data = 12'h3A7;
        15'h0073: data = 12'h0C4;
        15'h0074: data = 12'h766;
        15'h0075: data = 12'h5D5;
        15'h0076: data = 12'h04D;
        15'h0077: data = 12'h5B0;
        15'h0078: data = 12'h750;
        15'h0079: data = 12'h0AE;
        15'h007A: data = 12'h341;
        15'h007B: data = 12'h7F4;
        15'h007C: data = 12'h26D;
        15'h007D: data = 12'h172;
        15'h007E: data = 12'h7EC;
        15'h007F: data = 12'h474;
        15'h0080: data = 12'h08B;
        15'h0081: data = 12'h719;
        15'h0082: data = 12'h631;
        15'h0083: data = 12'h044;
        15'h0084: data = 12'h4BC;
        15'h0085: data = 12'h78C;
        15'h0086: data = 12'h146;
        15'h0087: data = 12'h271;
        15'h0088: data = 12'h805;
        15'h0089: data = 12'h357;
        15'h008A: data = 12'h7E7;
        15'h008B: data = 12'h7EB;
        15'h008C: data = 12'h7EC;
        15'h008D: data = 12'h7E7;
        15'h008E: data = 12'h7E9;
        15'h008F: data = 12'h7E9;
        15'h0090: data = 12'h7EA;
        15'h0091: data = 12'h7EC;
        15'h0092: data = 12'h7EA;
        15'h0093: data = 12'h7F2;
        15'h0094: data = 12'h7F6;
        15'h0095: data = 12'h7FA;
        15'h0096: data = 12'h7FC;
        15'h0097: data = 12'h7FE;
        15'h0098: data = 12'h7FE;
        15'h0099: data = 12'h800;
        15'h009A: data = 12'h7F7;
        15'h009B: data = 12'h7FA;
        15'h009C: data = 12'h7F9;
        15'h009D: data = 12'h7F8;
        15'h009E: data = 12'h7F6;
        15'h009F: data = 12'h7F5;
        15'h00A0: data = 12'h7F2;
        15'h00A1: data = 12'h7F0;
        15'h00A2: data = 12'h7F2;
        15'h00A3: data = 12'h7F4;
        15'h00A4: data = 12'h7FB;
        15'h00A5: data = 12'h802;
        15'h00A6: data = 12'h803;
        15'h00A7: data = 12'h805;
        15'h00A8: data = 12'h805;
        15'h00A9: data = 12'h803;
        15'h00AA: data = 12'h801;
        15'h00AB: data = 12'h7FB;
        15'h00AC: data = 12'h7FD;
        15'h00AD: data = 12'h7F9;
        15'h00AE: data = 12'h7F8;
        15'h00AF: data = 12'h7F8;
        15'h00B0: data = 12'h7F6;
        15'h00B1: data = 12'h7FE;
        15'h00B2: data = 12'h7FC;
        15'h00B3: data = 12'h801;
        15'h00B4: data = 12'h804;
        15'h00B5: data = 12'h805;
        15'h00B6: data = 12'h802;
        15'h00B7: data = 12'h803;
        15'h00B8: data = 12'h7F9;
        15'h00B9: data = 12'h7F9;
        15'h00BA: data = 12'h7F8;
        15'h00BB: data = 12'h7FA;
        15'h00BC: data = 12'h7FA;
        15'h00BD: data = 12'h7FD;
        15'h00BE: data = 12'h7FE;
        15'h00BF: data = 12'h807;
        15'h00C0: data = 12'h806;
        15'h00C1: data = 12'h805;
        15'h00C2: data = 12'h802;
        15'h00C3: data = 12'h7FD;
        15'h00C4: data = 12'h7FA;
        15'h00C5: data = 12'h7F7;
        15'h00C6: data = 12'h7F6;
        15'h00C7: data = 12'h7F8;
        15'h00C8: data = 12'h7FF;
        15'h00C9: data = 12'h801;
        15'h00CA: data = 12'h80A;
        15'h00CB: data = 12'h802;
        15'h00CC: data = 12'h804;
        15'h00CD: data = 12'h7FD;
        15'h00CE: data = 12'h7FB;
        15'h00CF: data = 12'h7F9;
        15'h00D0: data = 12'h7F5;
        15'h00D1: data = 12'h7FF;
        15'h00D2: data = 12'h801;
        15'h00D3: data = 12'h804;
        15'h00D4: data = 12'h804;
        15'h00D5: data = 12'h804;
        15'h00D6: data = 12'h7FF;
        15'h00D7: data = 12'h7FB;
        15'h00D8: data = 12'h7D8;
        15'h00D9: data = 12'h7DA;
        15'h00DA: data = 12'h7D8;
        15'h00DB: data = 12'h7E1;
        15'h00DC: data = 12'h7E2;
        15'h00DD: data = 12'h7DE;
        15'h00DE: data = 12'h7E3;
        15'h00DF: data = 12'h7E0;
        15'h00E0: data = 12'h7DB;
        15'h00E1: data = 12'h7D8;
        15'h00E2: data = 12'h7D8;
        15'h00E3: data = 12'h7DC;
        15'h00E4: data = 12'h7E2;
        15'h00E5: data = 12'h7E3;
        15'h00E6: data = 12'h7E3;
        15'h00E7: data = 12'h7E4;
        15'h00E8: data = 12'h7D9;
        15'h00E9: data = 12'h7D5;
        15'h00EA: data = 12'h7D2;
        15'h00EB: data = 12'h7D2;
        15'h00EC: data = 12'h7DC;
        15'h00ED: data = 12'h7DF;
        15'h00EE: data = 12'h7E6;
        15'h00EF: data = 12'h7E6;
        15'h00F0: data = 12'h7E2;
        15'h00F1: data = 12'h7DD;
        15'h00F2: data = 12'h7D6;
        15'h00F3: data = 12'h7D5;
        15'h00F4: data = 12'h7D5;
        15'h00F5: data = 12'h7D9;
        15'h00F6: data = 12'h7DE;
        15'h00F7: data = 12'h7E5;
        15'h00F8: data = 12'h7E3;
        15'h00F9: data = 12'h7E4;
        15'h00FA: data = 12'h7DC;
        15'h00FB: data = 12'h7D6;
        15'h00FC: data = 12'h7D1;
        15'h00FD: data = 12'h7D6;
        15'h00FE: data = 12'h7DB;
        15'h00FF: data = 12'h7E3;
        15'h0100: data = 12'h7E1;
        15'h0101: data = 12'h7E5;
        15'h0102: data = 12'h7E1;
        15'h0103: data = 12'h7D5;
        15'h0104: data = 12'h7D4;
        15'h0105: data = 12'h7D2;
        15'h0106: data = 12'h7D9;
        15'h0107: data = 12'h7E0;
        15'h0108: data = 12'h7E2;
        15'h0109: data = 12'h7E3;
        15'h010A: data = 12'h7E0;
        15'h010B: data = 12'h7DC;
        15'h010C: data = 12'h7D7;
        15'h010D: data = 12'h7D1;
        15'h010E: data = 12'h7D3;
        15'h010F: data = 12'h7D9;
        15'h0110: data = 12'h7DF;
        15'h0111: data = 12'h7E5;
        15'h0112: data = 12'h7E1;
        15'h0113: data = 12'h7DD;
        15'h0114: data = 12'h7D5;
        15'h0115: data = 12'h7D4;
        15'h0116: data = 12'h7D6;
        15'h0117: data = 12'h7DA;
        15'h0118: data = 12'h7DC;
        15'h0119: data = 12'h7DF;
        15'h011A: data = 12'h7C1;
        15'h011B: data = 12'h7C0;
        15'h011C: data = 12'h7BF;
        15'h011D: data = 12'h7B7;
        15'h011E: data = 12'h7B7;
        15'h011F: data = 12'h7B4;
        15'h0120: data = 12'h7BA;
        15'h0121: data = 12'h7BA;
        15'h0122: data = 12'h7C4;
        15'h0123: data = 12'h7C1;
        15'h0124: data = 12'h7C2;
        15'h0125: data = 12'h7BD;
        15'h0126: data = 12'h7B4;
        15'h0127: data = 12'h7B5;
        15'h0128: data = 12'h7B6;
        15'h0129: data = 12'h7B9;
        15'h012A: data = 12'h7BF;
        15'h012B: data = 12'h7C1;
        15'h012C: data = 12'h7C3;
        15'h012D: data = 12'h7C4;
        15'h012E: data = 12'h7BB;
        15'h012F: data = 12'h7BB;
        15'h0130: data = 12'h7B7;
        15'h0131: data = 12'h7B4;
        15'h0132: data = 12'h7B9;
        15'h0133: data = 12'h7BB;
        15'h0134: data = 12'h7C2;
        15'h0135: data = 12'h7BF;
        15'h0136: data = 12'h7BB;
        15'h0137: data = 12'h7BC;
        15'h0138: data = 12'h7B5;
        15'h0139: data = 12'h7B1;
        15'h013A: data = 12'h7B5;
        15'h013B: data = 12'h7B6;
        15'h013C: data = 12'h7BD;
        15'h013D: data = 12'h7C0;
        15'h013E: data = 12'h7C0;
        15'h013F: data = 12'h7C1;
        15'h0140: data = 12'h7BB;
        15'h0141: data = 12'h7B8;
        15'h0142: data = 12'h7B6;
        15'h0143: data = 12'h7B7;
        15'h0144: data = 12'h7B3;
        15'h0145: data = 12'h7BE;
        15'h0146: data = 12'h7BF;
        15'h0147: data = 12'h7C1;
        15'h0148: data = 12'h7C1;
        15'h0149: data = 12'h7C3;
        15'h014A: data = 12'h7BE;
        15'h014B: data = 12'h7BB;
        15'h014C: data = 12'h7B5;
        15'h014D: data = 12'h7B8;
        15'h014E: data = 12'h7B8;
        15'h014F: data = 12'h7BB;
        15'h0150: data = 12'h7BB;
        15'h0151: data = 12'h7C0;
        15'h0152: data = 12'h7C0;
        15'h0153: data = 12'h7BF;
        15'h0154: data = 12'h7B6;
        15'h0155: data = 12'h7B9;
        15'h0156: data = 12'h7B5;
        15'h0157: data = 12'h7B3;
        15'h0158: data = 12'h7B8;
        15'h0159: data = 12'h7BA;
        15'h015A: data = 12'h7BF;
        15'h015B: data = 12'h7C0;
        15'h015C: data = 12'h7BC;
        15'h015D: data = 12'h7BE;
        15'h015E: data = 12'h7B8;
        15'h015F: data = 12'h7B6;
        15'h0160: data = 12'h7B6;
        15'h0161: data = 12'h7B7;
        15'h0162: data = 12'h7B7;
        15'h0163: data = 12'h7BA;
        15'h0164: data = 12'h7BC;
        15'h0165: data = 12'h7BD;
        15'h0166: data = 12'h7BC;
        15'h0167: data = 12'h7B8;
        15'h0168: data = 12'h797;
        15'h0169: data = 12'h795;
        15'h016A: data = 12'h797;
        15'h016B: data = 12'h795;
        15'h016C: data = 12'h794;
        15'h016D: data = 12'h79D;
        15'h016E: data = 12'h79D;
        15'h016F: data = 12'h7A2;
        15'h0170: data = 12'h7A1;
        15'h0171: data = 12'h79E;
        15'h0172: data = 12'h79A;
        15'h0173: data = 12'h792;
        15'h0174: data = 12'h792;
        15'h0175: data = 12'h795;
        15'h0176: data = 12'h797;
        15'h0177: data = 12'h79A;
        15'h0178: data = 12'h79B;
        15'h0179: data = 12'h7A4;
        15'h017A: data = 12'h79D;
        15'h017B: data = 12'h799;
        15'h017C: data = 12'h796;
        15'h017D: data = 12'h797;
        15'h017E: data = 12'h797;
        15'h017F: data = 12'h791;
        15'h0180: data = 12'h79B;
        15'h0181: data = 12'h79E;
        15'h0182: data = 12'h79F;
        15'h0183: data = 12'h7A4;
        15'h0184: data = 12'h79F;
        15'h0185: data = 12'h79F;
        15'h0186: data = 12'h799;
        15'h0187: data = 12'h793;
        15'h0188: data = 12'h793;
        15'h0189: data = 12'h794;
        15'h018A: data = 12'h798;
        15'h018B: data = 12'h79F;
        15'h018C: data = 12'h79D;
        15'h018D: data = 12'h7A0;
        15'h018E: data = 12'h79D;
        15'h018F: data = 12'h799;
        15'h0190: data = 12'h799;
        15'h0191: data = 12'h790;
        15'h0192: data = 12'h793;
        15'h0193: data = 12'h794;
        15'h0194: data = 12'h797;
        15'h0195: data = 12'h7A3;
        15'h0196: data = 12'h7A3;
        15'h0197: data = 12'h79E;
        15'h0198: data = 12'h7A1;
        15'h0199: data = 12'h79A;
        15'h019A: data = 12'h797;
        15'h019B: data = 12'h793;
        15'h019C: data = 12'h78F;
        15'h019D: data = 12'h796;
        15'h019E: data = 12'h798;
        15'h019F: data = 12'h79D;
        15'h01A0: data = 12'h7A3;
        15'h01A1: data = 12'h7A2;
        15'h01A2: data = 12'h7A0;
        15'h01A3: data = 12'h79D;
        15'h01A4: data = 12'h798;
        15'h01A5: data = 12'h796;
        15'h01A6: data = 12'h796;
        15'h01A7: data = 12'h79A;
        15'h01A8: data = 12'h79D;
        15'h01A9: data = 12'h79E;
        15'h01AA: data = 12'h780;
        15'h01AB: data = 12'h77F;
        15'h01AC: data = 12'h77D;
        15'h01AD: data = 12'h779;
        15'h01AE: data = 12'h775;
        15'h01AF: data = 12'h774;
        15'h01B0: data = 12'h778;
        15'h01B1: data = 12'h77D;
        15'h01B2: data = 12'h77D;
        15'h01B3: data = 12'h781;
        15'h01B4: data = 12'h781;
        15'h01B5: data = 12'h780;
        15'h01B6: data = 12'h77B;
        15'h01B7: data = 12'h779;
        15'h01B8: data = 12'h775;
        15'h01B9: data = 12'h776;
        15'h01BA: data = 12'h778;
        15'h01BB: data = 12'h77F;
        default: data = 12'h000;
    endcase
end

endmodule

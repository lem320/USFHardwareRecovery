module rom_test (
    input [14:0] address,
    output reg [11:0] data
);

always @(*) begin
    case (address)
        15'h0000: data = 12'h349;
        15'h0001: data = 12'h34B;
        15'h0002: data = 12'h350;
        15'h0003: data = 12'h354;
        15'h0004: data = 12'h355;
        15'h0005: data = 12'h355;
        15'h0006: data = 12'h354;
        15'h0007: data = 12'h34E;
        15'h0008: data = 12'h34E;
        15'h0009: data = 12'h348;
        15'h000A: data = 12'h34C;
        15'h000B: data = 12'h34D;
        15'h000C: data = 12'h34F;
        15'h000D: data = 12'h354;
        15'h000E: data = 12'h353;
        15'h000F: data = 12'h355;
        15'h0010: data = 12'h353;
        15'h0011: data = 12'h351;
        15'h0012: data = 12'h34C;
        15'h0013: data = 12'h34A;
        15'h0014: data = 12'h349;
        15'h0015: data = 12'h34C;
        15'h0016: data = 12'h351;
        15'h0017: data = 12'h354;
        15'h0018: data = 12'h353;
        15'h0019: data = 12'h350;
        15'h001A: data = 12'h34A;
        15'h001B: data = 12'h349;
        15'h001C: data = 12'h349;
        15'h001D: data = 12'h349;
        15'h001E: data = 12'h34C;
        15'h001F: data = 12'h355;
        15'h0020: data = 12'h353;
        15'h0021: data = 12'h351;
        15'h0022: data = 12'h34F;
        15'h0023: data = 12'h34C;
        15'h0024: data = 12'h34D;
        15'h0025: data = 12'h34A;
        15'h0026: data = 12'h351;
        15'h0027: data = 12'h352;
        15'h0028: data = 12'h355;
        15'h0029: data = 12'h354;
        15'h002A: data = 12'h356;
        15'h002B: data = 12'h351;
        15'h002C: data = 12'h34B;
        15'h002D: data = 12'h346;
        15'h002E: data = 12'h346;
        15'h002F: data = 12'h346;
        15'h0030: data = 12'h34F;
        15'h0031: data = 12'h354;
        15'h0032: data = 12'h355;
        15'h0033: data = 12'h358;
        15'h0034: data = 12'h353;
        15'h0035: data = 12'h34F;
        15'h0036: data = 12'h34A;
        15'h0037: data = 12'h348;
        15'h0038: data = 12'h34C;
        15'h0039: data = 12'h34B;
        15'h003A: data = 12'h351;
        15'h003B: data = 12'h356;
        15'h003C: data = 12'h356;
        15'h003D: data = 12'h355;
        15'h003E: data = 12'h34E;
        15'h003F: data = 12'h34C;
        15'h0040: data = 12'h34A;
        15'h0041: data = 12'h347;
        15'h0042: data = 12'h34D;
        15'h0043: data = 12'h352;
        15'h0044: data = 12'h354;
        15'h0045: data = 12'h357;
        15'h0046: data = 12'h358;
        15'h0047: data = 12'h34F;
        15'h0048: data = 12'h34C;
        15'h0049: data = 12'h349;
        15'h004A: data = 12'h343;
        15'h004B: data = 12'h345;
        15'h004C: data = 12'h34F;
        15'h004D: data = 12'h357;
        15'h004E: data = 12'h353;
        15'h004F: data = 12'h356;
        15'h0050: data = 12'h352;
        15'h0051: data = 12'h34F;
        15'h0052: data = 12'h348;
        15'h0053: data = 12'h349;
        15'h0054: data = 12'h34B;
        15'h0055: data = 12'h34D;
        15'h0056: data = 12'h352;
        15'h0057: data = 12'h355;
        15'h0058: data = 12'h354;
        15'h0059: data = 12'h356;
        15'h005A: data = 12'h351;
        15'h005B: data = 12'h34B;
        15'h005C: data = 12'h349;
        15'h005D: data = 12'h34B;
        15'h005E: data = 12'h34A;
        15'h005F: data = 12'h351;
        15'h0060: data = 12'h375;
        15'h0061: data = 12'h37B;
        15'h0062: data = 12'h375;
        15'h0063: data = 12'h373;
        15'h0064: data = 12'h370;
        15'h0065: data = 12'h36E;
        15'h0066: data = 12'h36A;
        15'h0067: data = 12'h36C;
        15'h0068: data = 12'h371;
        15'h0069: data = 12'h375;
        15'h006A: data = 12'h375;
        15'h006B: data = 12'h377;
        15'h006C: data = 12'h375;
        15'h006D: data = 12'h373;
        15'h006E: data = 12'h36B;
        15'h006F: data = 12'h36A;
        15'h0070: data = 12'h36C;
        15'h0071: data = 12'h36C;
        15'h0072: data = 12'h370;
        15'h0073: data = 12'h373;
        15'h0074: data = 12'h374;
        15'h0075: data = 12'h372;
        15'h0076: data = 12'h373;
        15'h0077: data = 12'h36B;
        15'h0078: data = 12'h36B;
        15'h0079: data = 12'h36B;
        15'h007A: data = 12'h36A;
        15'h007B: data = 12'h36E;
        15'h007C: data = 12'h373;
        15'h007D: data = 12'h379;
        15'h007E: data = 12'h375;
        15'h007F: data = 12'h371;
        15'h0080: data = 12'h371;
        15'h0081: data = 12'h369;
        15'h0082: data = 12'h36A;
        15'h0083: data = 12'h36D;
        15'h0084: data = 12'h36D;
        15'h0085: data = 12'h375;
        15'h0086: data = 12'h378;
        15'h0087: data = 12'h378;
        15'h0088: data = 12'h376;
        15'h0089: data = 12'h372;
        15'h008A: data = 12'h36C;
        15'h008B: data = 12'h36D;
        15'h008C: data = 12'h368;
        15'h008D: data = 12'h36F;
        15'h008E: data = 12'h376;
        15'h008F: data = 12'h378;
        15'h0090: data = 12'h374;
        15'h0091: data = 12'h37A;
        15'h0092: data = 12'h373;
        15'h0093: data = 12'h36C;
        15'h0094: data = 12'h369;
        15'h0095: data = 12'h369;
        15'h0096: data = 12'h36C;
        15'h0097: data = 12'h36F;
        15'h0098: data = 12'h375;
        15'h0099: data = 12'h376;
        15'h009A: data = 12'h378;
        15'h009B: data = 12'h375;
        15'h009C: data = 12'h373;
        15'h009D: data = 12'h36A;
        15'h009E: data = 12'h36A;
        15'h009F: data = 12'h367;
        15'h00A0: data = 12'h36D;
        15'h00A1: data = 12'h373;
        15'h00A2: data = 12'h376;
        15'h00A3: data = 12'h37A;
        15'h00A4: data = 12'h373;
        15'h00A5: data = 12'h371;
        15'h00A6: data = 12'h36B;
        15'h00A7: data = 12'h368;
        15'h00A8: data = 12'h368;
        15'h00A9: data = 12'h36F;
        15'h00AA: data = 12'h371;
        15'h00AB: data = 12'h377;
        15'h00AC: data = 12'h372;
        15'h00AD: data = 12'h372;
        15'h00AE: data = 12'h36F;
        15'h00AF: data = 12'h36A;
        15'h00B0: data = 12'h366;
        15'h00B1: data = 12'h368;
        15'h00B2: data = 12'h36A;
        15'h00B3: data = 12'h36F;
        15'h00B4: data = 12'h374;
        15'h00B5: data = 12'h375;
        15'h00B6: data = 12'h372;
        15'h00B7: data = 12'h374;
        15'h00B8: data = 12'h36C;
        15'h00B9: data = 12'h36A;
        15'h00BA: data = 12'h368;
        15'h00BB: data = 12'h36A;
        15'h00BC: data = 12'h38B;
        15'h00BD: data = 12'h38B;
        15'h00BE: data = 12'h391;
        15'h00BF: data = 12'h390;
        15'h00C0: data = 12'h392;
        15'h00C1: data = 12'h395;
        15'h00C2: data = 12'h390;
        15'h00C3: data = 12'h388;
        15'h00C4: data = 12'h389;
        15'h00C5: data = 12'h387;
        15'h00C6: data = 12'h38C;
        15'h00C7: data = 12'h391;
        15'h00C8: data = 12'h397;
        15'h00C9: data = 12'h399;
        15'h00CA: data = 12'h396;
        15'h00CB: data = 12'h38E;
        15'h00CC: data = 12'h388;
        15'h00CD: data = 12'h389;
        15'h00CE: data = 12'h387;
        15'h00CF: data = 12'h38B;
        15'h00D0: data = 12'h396;
        15'h00D1: data = 12'h397;
        15'h00D2: data = 12'h397;
        15'h00D3: data = 12'h397;
        15'h00D4: data = 12'h38E;
        15'h00D5: data = 12'h38A;
        15'h00D6: data = 12'h388;
        15'h00D7: data = 12'h389;
        15'h00D8: data = 12'h38F;
        15'h00D9: data = 12'h392;
        15'h00DA: data = 12'h397;
        15'h00DB: data = 12'h394;
        15'h00DC: data = 12'h394;
        15'h00DD: data = 12'h391;
        15'h00DE: data = 12'h38B;
        15'h00DF: data = 12'h387;
        15'h00E0: data = 12'h38B;
        15'h00E1: data = 12'h38A;
        15'h00E2: data = 12'h392;
        15'h00E3: data = 12'h394;
        15'h00E4: data = 12'h397;
        15'h00E5: data = 12'h394;
        15'h00E6: data = 12'h391;
        15'h00E7: data = 12'h38E;
        15'h00E8: data = 12'h388;
        15'h00E9: data = 12'h388;
        15'h00EA: data = 12'h386;
        15'h00EB: data = 12'h38D;
        15'h00EC: data = 12'h396;
        15'h00ED: data = 12'h396;
        15'h00EE: data = 12'h397;
        15'h00EF: data = 12'h393;
        15'h00F0: data = 12'h38E;
        15'h00F1: data = 12'h388;
        15'h00F2: data = 12'h386;
        15'h00F3: data = 12'h389;
        15'h00F4: data = 12'h38A;
        15'h00F5: data = 12'h392;
        15'h00F6: data = 12'h396;
        15'h00F7: data = 12'h399;
        15'h00F8: data = 12'h398;
        15'h00F9: data = 12'h392;
        15'h00FA: data = 12'h38F;
        15'h00FB: data = 12'h387;
        15'h00FC: data = 12'h387;
        15'h00FD: data = 12'h38B;
        15'h00FE: data = 12'h38D;
        15'h00FF: data = 12'h398;
        15'h0100: data = 12'h396;
        15'h0101: data = 12'h397;
        15'h0102: data = 12'h390;
        15'h0103: data = 12'h38B;
        15'h0104: data = 12'h38B;
        15'h0105: data = 12'h387;
        15'h0106: data = 12'h38C;
        15'h0107: data = 12'h389;
        15'h0108: data = 12'h392;
        15'h0109: data = 12'h395;
        15'h010A: data = 12'h393;
        15'h010B: data = 12'h395;
        15'h010C: data = 12'h391;
        15'h010D: data = 12'h38B;
        15'h010E: data = 12'h38A;
        15'h010F: data = 12'h388;
        15'h0110: data = 12'h389;
        15'h0111: data = 12'h38C;
        15'h0112: data = 12'h390;
        15'h0113: data = 12'h395;
        15'h0114: data = 12'h395;
        15'h0115: data = 12'h396;
        15'h0116: data = 12'h38C;
        15'h0117: data = 12'h39B;
        15'h0118: data = 12'h3A8;
        15'h0119: data = 12'h3A9;
        15'h011A: data = 12'h3AC;
        15'h011B: data = 12'h3B2;
        15'h011C: data = 12'h3B5;
        15'h011D: data = 12'h3B7;
        15'h011E: data = 12'h3B8;
        15'h011F: data = 12'h3AE;
        15'h0120: data = 12'h3AA;
        15'h0121: data = 12'h3AB;
        15'h0122: data = 12'h3A6;
        15'h0123: data = 12'h3AA;
        15'h0124: data = 12'h3AE;
        15'h0125: data = 12'h3B1;
        15'h0126: data = 12'h3B5;
        15'h0127: data = 12'h3B2;
        15'h0128: data = 12'h3AF;
        15'h0129: data = 12'h3AA;
        15'h012A: data = 12'h3A9;
        15'h012B: data = 12'h3AA;
        15'h012C: data = 12'h3AB;
        15'h012D: data = 12'h3B2;
        15'h012E: data = 12'h3B6;
        15'h012F: data = 12'h3B3;
        15'h0130: data = 12'h3B5;
        15'h0131: data = 12'h3B0;
        15'h0132: data = 12'h3AF;
        15'h0133: data = 12'h3A8;
        15'h0134: data = 12'h3A5;
        15'h0135: data = 12'h3A7;
        15'h0136: data = 12'h3AF;
        15'h0137: data = 12'h3B1;
        15'h0138: data = 12'h3B5;
        15'h0139: data = 12'h3B5;
        15'h013A: data = 12'h3B1;
        15'h013B: data = 12'h3AD;
        15'h013C: data = 12'h3AA;
        15'h013D: data = 12'h3A7;
        15'h013E: data = 12'h3AC;
        15'h013F: data = 12'h3AA;
        15'h0140: data = 12'h3B0;
        15'h0141: data = 12'h3B6;
        15'h0142: data = 12'h3B6;
        15'h0143: data = 12'h3B1;
        15'h0144: data = 12'h3B0;
        15'h0145: data = 12'h3AC;
        15'h0146: data = 12'h3A7;
        15'h0147: data = 12'h3A6;
        15'h0148: data = 12'h3AA;
        15'h0149: data = 12'h3AE;
        15'h014A: data = 12'h3B2;
        15'h014B: data = 12'h3B6;
        15'h014C: data = 12'h3B4;
        15'h014D: data = 12'h3B3;
        15'h014E: data = 12'h3AC;
        15'h014F: data = 12'h3AB;
        15'h0150: data = 12'h3AA;
        15'h0151: data = 12'h3A8;
        15'h0152: data = 12'h3AE;
        15'h0153: data = 12'h3B2;
        15'h0154: data = 12'h3B3;
        15'h0155: data = 12'h3B4;
        15'h0156: data = 12'h3B5;
        15'h0157: data = 12'h3AF;
        15'h0158: data = 12'h3AB;
        15'h0159: data = 12'h3A8;
        15'h015A: data = 12'h3A7;
        15'h015B: data = 12'h3AA;
        15'h015C: data = 12'h3B0;
        15'h015D: data = 12'h3B6;
        15'h015E: data = 12'h3B4;
        15'h015F: data = 12'h3B1;
        15'h0160: data = 12'h3B4;
        15'h0161: data = 12'h3AC;
        15'h0162: data = 12'h3A9;
        15'h0163: data = 12'h3AA;
        15'h0164: data = 12'h3A9;
        15'h0165: data = 12'h3B2;
        15'h0166: data = 12'h3B5;
        15'h0167: data = 12'h3BA;
        15'h0168: data = 12'h3BA;
        15'h0169: data = 12'h3B3;
        15'h016A: data = 12'h3AD;
        15'h016B: data = 12'h3A9;
        15'h016C: data = 12'h3A6;
        15'h016D: data = 12'h3A7;
        15'h016E: data = 12'h3AE;
        15'h016F: data = 12'h3B2;
        15'h0170: data = 12'h3B8;
        15'h0171: data = 12'h3B4;
        15'h0172: data = 12'h3B0;
        15'h0173: data = 12'h3AE;
        15'h0174: data = 12'h3A9;
        15'h0175: data = 12'h3A4;
        15'h0176: data = 12'h3A9;
        15'h0177: data = 12'h3AE;
        15'h0178: data = 12'h3B1;
        15'h0179: data = 12'h3B8;
        15'h017A: data = 12'h3B7;
        15'h017B: data = 12'h3B3;
        15'h017C: data = 12'h3AF;
        15'h017D: data = 12'h3A9;
        15'h017E: data = 12'h3A9;
        15'h017F: data = 12'h3A8;
        15'h0180: data = 12'h3CE;
        15'h0181: data = 12'h3D1;
        15'h0182: data = 12'h3D7;
        15'h0183: data = 12'h3D6;
        15'h0184: data = 12'h3D1;
        15'h0185: data = 12'h3D2;
        15'h0186: data = 12'h3CF;
        15'h0187: data = 12'h3CB;
        15'h0188: data = 12'h3C6;
        15'h0189: data = 12'h3CA;
        15'h018A: data = 12'h3D0;
        15'h018B: data = 12'h3D3;
        15'h018C: data = 12'h3D3;
        15'h018D: data = 12'h3D4;
        15'h018E: data = 12'h3D3;
        15'h018F: data = 12'h3CD;
        15'h0190: data = 12'h3C8;
        15'h0191: data = 12'h3C6;
        15'h0192: data = 12'h3C8;
        15'h0193: data = 12'h3CD;
        15'h0194: data = 12'h3D6;
        15'h0195: data = 12'h3D5;
        15'h0196: data = 12'h3D4;
        15'h0197: data = 12'h3D3;
        15'h0198: data = 12'h3CD;
        15'h0199: data = 12'h3CC;
        15'h019A: data = 12'h3CC;
        15'h019B: data = 12'h3C6;
        15'h019C: data = 12'h3CA;
        15'h019D: data = 12'h3D3;
        15'h019E: data = 12'h3D5;
        15'h019F: data = 12'h3D2;
        15'h01A0: data = 12'h3D1;
        15'h01A1: data = 12'h3D1;
        15'h01A2: data = 12'h3CC;
        15'h01A3: data = 12'h3CA;
        15'h01A4: data = 12'h3C5;
        15'h01A5: data = 12'h3C9;
        15'h01A6: data = 12'h3D0;
        15'h01A7: data = 12'h3D4;
        15'h01A8: data = 12'h3D6;
        15'h01A9: data = 12'h3D8;
        15'h01AA: data = 12'h3D6;
        15'h01AB: data = 12'h3CE;
        15'h01AC: data = 12'h3CC;
        15'h01AD: data = 12'h3C4;
        15'h01AE: data = 12'h3CA;
        15'h01AF: data = 12'h3CD;
        15'h01B0: data = 12'h3D1;
        15'h01B1: data = 12'h3D5;
        15'h01B2: data = 12'h3D3;
        15'h01B3: data = 12'h3D5;
        15'h01B4: data = 12'h3CC;
        15'h01B5: data = 12'h3CA;
        15'h01B6: data = 12'h3C8;
        15'h01B7: data = 12'h3C8;
        15'h01B8: data = 12'h3CE;
        15'h01B9: data = 12'h3D0;
        15'h01BA: data = 12'h3D5;
        15'h01BB: data = 12'h3D2;
        15'h01BC: data = 12'h3D3;
        15'h01BD: data = 12'h3CF;
        15'h01BE: data = 12'h3CB;
        15'h01BF: data = 12'h3CB;
        15'h01C0: data = 12'h3C8;
        15'h01C1: data = 12'h3CC;
        15'h01C2: data = 12'h3D5;
        15'h01C3: data = 12'h3D8;
        15'h01C4: data = 12'h3D6;
        15'h01C5: data = 12'h3D4;
        15'h01C6: data = 12'h3D3;
        15'h01C7: data = 12'h3CD;
        15'h01C8: data = 12'h3CB;
        15'h01C9: data = 12'h3CA;
        15'h01CA: data = 12'h3CB;
        15'h01CB: data = 12'h3CF;
        15'h01CC: data = 12'h3CF;
        15'h01CD: data = 12'h3D5;
        15'h01CE: data = 12'h3D3;
        15'h01CF: data = 12'h3D3;
        15'h01D0: data = 12'h3CE;
        15'h01D1: data = 12'h3CA;
        15'h01D2: data = 12'h3C6;
        15'h01D3: data = 12'h3CB;
        15'h01D4: data = 12'h3CD;
        15'h01D5: data = 12'h3D0;
        15'h01D6: data = 12'h3D7;
        15'h01D7: data = 12'h3D6;
        15'h01D8: data = 12'h3D4;
        15'h01D9: data = 12'h3CF;
        15'h01DA: data = 12'h3CC;
        15'h01DB: data = 12'h3C8;
        15'h01DC: data = 12'h3EB;
        15'h01DD: data = 12'h3EA;
        15'h01DE: data = 12'h3F1;
        15'h01DF: data = 12'h3F4;
        15'h01E0: data = 12'h3F7;
        15'h01E1: data = 12'h3F6;
        15'h01E2: data = 12'h3F3;
        15'h01E3: data = 12'h3EB;
        15'h01E4: data = 12'h3E7;
        15'h01E5: data = 12'h3EB;
        15'h01E6: data = 12'h3EB;
        15'h01E7: data = 12'h3EF;
        15'h01E8: data = 12'h3F5;
        15'h01E9: data = 12'h3FA;
        15'h01EA: data = 12'h3F5;
        15'h01EB: data = 12'h3F4;
        15'h01EC: data = 12'h3EE;
        15'h01ED: data = 12'h3EA;
        15'h01EE: data = 12'h3EB;
        15'h01EF: data = 12'h3EB;
        15'h01F0: data = 12'h3F3;
        15'h01F1: data = 12'h3F5;
        15'h01F2: data = 12'h3F5;
        15'h01F3: data = 12'h3F5;
        15'h01F4: data = 12'h3F1;
        15'h01F5: data = 12'h3EC;
        15'h01F6: data = 12'h3ED;
        15'h01F7: data = 12'h3E9;
        15'h01F8: data = 12'h3ED;
        15'h01F9: data = 12'h3EE;
        15'h01FA: data = 12'h3F3;
        15'h01FB: data = 12'h3F4;
        15'h01FC: data = 12'h3F5;
        15'h01FD: data = 12'h3F1;
        15'h01FE: data = 12'h3F2;
        15'h01FF: data = 12'h3EC;
        15'h0200: data = 12'h3EA;
        15'h0201: data = 12'h3ED;
        15'h0202: data = 12'h3EF;
        15'h0203: data = 12'h3EF;
        15'h0204: data = 12'h3F4;
        15'h0205: data = 12'h3F5;
        15'h0206: data = 12'h3F4;
        15'h0207: data = 12'h3F2;
        15'h0208: data = 12'h3EB;
        15'h0209: data = 12'h3ED;
        15'h020A: data = 12'h3E8;
        15'h020B: data = 12'h3E8;
        15'h020C: data = 12'h3F2;
        15'h020D: data = 12'h3F2;
        15'h020E: data = 12'h3F4;
        15'h020F: data = 12'h3F5;
        15'h0210: data = 12'h3F4;
        15'h0211: data = 12'h3EF;
        15'h0212: data = 12'h3ED;
        15'h0213: data = 12'h3EA;
        15'h0214: data = 12'h3EA;
        15'h0215: data = 12'h3EB;
        15'h0216: data = 12'h3F3;
        15'h0217: data = 12'h3F5;
        15'h0218: data = 12'h3F5;
        15'h0219: data = 12'h3F3;
        15'h021A: data = 12'h3F2;
        15'h021B: data = 12'h3EB;
        15'h021C: data = 12'h3EA;
        15'h021D: data = 12'h3E9;
        15'h021E: data = 12'h3ED;
        15'h021F: data = 12'h3F0;
        15'h0220: data = 12'h3F5;
        15'h0221: data = 12'h3F9;
        15'h0222: data = 12'h3F9;
        15'h0223: data = 12'h3F4;
        15'h0224: data = 12'h3EC;
        15'h0225: data = 12'h3EA;
        15'h0226: data = 12'h3E9;
        15'h0227: data = 12'h3ED;
        15'h0228: data = 12'h3F3;
        15'h0229: data = 12'h3F7;
        15'h022A: data = 12'h3F8;
        15'h022B: data = 12'h3F6;
        15'h022C: data = 12'h3F6;
        15'h022D: data = 12'h3F0;
        15'h022E: data = 12'h3EB;
        15'h022F: data = 12'h3E8;
        15'h0230: data = 12'h3F0;
        15'h0231: data = 12'h3F1;
        15'h0232: data = 12'h3F6;
        15'h0233: data = 12'h3FD;
        15'h0234: data = 12'h3F9;
        15'h0235: data = 12'h3F5;
        15'h0236: data = 12'h3F0;
        15'h0237: data = 12'h3ED;
        15'h0238: data = 12'h3EB;
        15'h0239: data = 12'h3EE;
        15'h023A: data = 12'h3F0;
        15'h023B: data = 12'h3F1;
        15'h023C: data = 12'h3F5;
        15'h023D: data = 12'h3F7;
        15'h023E: data = 12'h3F6;
        15'h023F: data = 12'h3F5;
        15'h0240: data = 12'h3ED;
        15'h0241: data = 12'h3E7;
        15'h0242: data = 12'h3E8;
        15'h0243: data = 12'h3EB;
        15'h0244: data = 12'h3EF;
        15'h0245: data = 12'h416;
        15'h0246: data = 12'h419;
        15'h0247: data = 12'h419;
        15'h0248: data = 12'h417;
        15'h0249: data = 12'h40D;
        15'h024A: data = 12'h40C;
        15'h024B: data = 12'h409;
        15'h024C: data = 12'h40A;
        15'h024D: data = 12'h410;
        15'h024E: data = 12'h418;
        15'h024F: data = 12'h414;
        15'h0250: data = 12'h418;
        15'h0251: data = 12'h412;
        15'h0252: data = 12'h411;
        15'h0253: data = 12'h409;
        15'h0254: data = 12'h408;
        15'h0255: data = 12'h40D;
        15'h0256: data = 12'h40D;
        15'h0257: data = 12'h414;
        15'h0258: data = 12'h414;
        15'h0259: data = 12'h416;
        15'h025A: data = 12'h413;
        15'h025B: data = 12'h411;
        15'h025C: data = 12'h40D;
        15'h025D: data = 12'h40B;
        15'h025E: data = 12'h40B;
        15'h025F: data = 12'h40B;
        15'h0260: data = 12'h413;
        15'h0261: data = 12'h414;
        15'h0262: data = 12'h412;
        15'h0263: data = 12'h419;
        15'h0264: data = 12'h414;
        15'h0265: data = 12'h40E;
        15'h0266: data = 12'h40A;
        15'h0267: data = 12'h40A;
        15'h0268: data = 12'h405;
        15'h0269: data = 12'h40F;
        15'h026A: data = 12'h414;
        15'h026B: data = 12'h416;
        15'h026C: data = 12'h418;
        15'h026D: data = 12'h415;
        15'h026E: data = 12'h411;
        15'h026F: data = 12'h40C;
        15'h0270: data = 12'h409;
        15'h0271: data = 12'h405;
        15'h0272: data = 12'h40B;
        15'h0273: data = 12'h413;
        15'h0274: data = 12'h417;
        15'h0275: data = 12'h418;
        15'h0276: data = 12'h414;
        15'h0277: data = 12'h40A;
        15'h0278: data = 12'h405;
        15'h0279: data = 12'h409;
        15'h027A: data = 12'h40A;
        15'h027B: data = 12'h40A;
        15'h027C: data = 12'h412;
        15'h027D: data = 12'h415;
        15'h027E: data = 12'h41A;
        15'h027F: data = 12'h417;
        15'h0280: data = 12'h413;
        15'h0281: data = 12'h40E;
        15'h0282: data = 12'h408;
        15'h0283: data = 12'h40C;
        15'h0284: data = 12'h40A;
        15'h0285: data = 12'h40E;
        15'h0286: data = 12'h418;
        15'h0287: data = 12'h419;
        15'h0288: data = 12'h41B;
        15'h0289: data = 12'h417;
        15'h028A: data = 12'h410;
        15'h028B: data = 12'h407;
        15'h028C: data = 12'h408;
        15'h028D: data = 12'h40B;
        15'h028E: data = 12'h413;
        15'h028F: data = 12'h41B;
        15'h0290: data = 12'h41C;
        15'h0291: data = 12'h419;
        15'h0292: data = 12'h410;
        15'h0293: data = 12'h40C;
        15'h0294: data = 12'h408;
        15'h0295: data = 12'h408;
        15'h0296: data = 12'h40C;
        15'h0297: data = 12'h412;
        15'h0298: data = 12'h416;
        15'h0299: data = 12'h418;
        15'h029A: data = 12'h416;
        15'h029B: data = 12'h415;
        15'h029C: data = 12'h410;
        15'h029D: data = 12'h407;
        15'h029E: data = 12'h40B;
        15'h029F: data = 12'h40E;
        15'h02A0: data = 12'h40F;
        15'h02A1: data = 12'h435;
        15'h02A2: data = 12'h436;
        15'h02A3: data = 12'h433;
        15'h02A4: data = 12'h436;
        15'h02A5: data = 12'h432;
        15'h02A6: data = 12'h42F;
        15'h02A7: data = 12'h42C;
        15'h02A8: data = 12'h42C;
        15'h02A9: data = 12'h429;
        15'h02AA: data = 12'h432;
        15'h02AB: data = 12'h431;
        15'h02AC: data = 12'h434;
        15'h02AD: data = 12'h435;
        15'h02AE: data = 12'h433;
        15'h02AF: data = 12'h434;
        15'h02B0: data = 12'h42D;
        15'h02B1: data = 12'h428;
        15'h02B2: data = 12'h42B;
        15'h02B3: data = 12'h42E;
        15'h02B4: data = 12'h42F;
        15'h02B5: data = 12'h434;
        15'h02B6: data = 12'h433;
        15'h02B7: data = 12'h432;
        15'h02B8: data = 12'h42C;
        15'h02B9: data = 12'h42B;
        15'h02BA: data = 12'h425;
        15'h02BB: data = 12'h426;
        15'h02BC: data = 12'h42C;
        15'h02BD: data = 12'h434;
        15'h02BE: data = 12'h433;
        15'h02BF: data = 12'h435;
        15'h02C0: data = 12'h431;
        15'h02C1: data = 12'h430;
        15'h02C2: data = 12'h42C;
        15'h02C3: data = 12'h427;
        15'h02C4: data = 12'h42C;
        15'h02C5: data = 12'h42E;
        15'h02C6: data = 12'h430;
        15'h02C7: data = 12'h432;
        15'h02C8: data = 12'h436;
        15'h02C9: data = 12'h434;
        15'h02CA: data = 12'h431;
        15'h02CB: data = 12'h42D;
        15'h02CC: data = 12'h42B;
        15'h02CD: data = 12'h426;
        15'h02CE: data = 12'h42B;
        15'h02CF: data = 12'h42C;
        15'h02D0: data = 12'h434;
        15'h02D1: data = 12'h438;
        15'h02D2: data = 12'h438;
        15'h02D3: data = 12'h433;
        15'h02D4: data = 12'h430;
        15'h02D5: data = 12'h42A;
        15'h02D6: data = 12'h427;
        15'h02D7: data = 12'h42B;
        15'h02D8: data = 12'h42E;
        15'h02D9: data = 12'h432;
        15'h02DA: data = 12'h437;
        15'h02DB: data = 12'h436;
        15'h02DC: data = 12'h434;
        15'h02DD: data = 12'h430;
        15'h02DE: data = 12'h429;
        15'h02DF: data = 12'h428;
        15'h02E0: data = 12'h428;
        15'h02E1: data = 12'h42C;
        15'h02E2: data = 12'h433;
        15'h02E3: data = 12'h435;
        15'h02E4: data = 12'h43A;
        15'h02E5: data = 12'h438;
        15'h02E6: data = 12'h433;
        15'h02E7: data = 12'h42B;
        15'h02E8: data = 12'h428;
        15'h02E9: data = 12'h428;
        15'h02EA: data = 12'h42C;
        15'h02EB: data = 12'h42E;
        15'h02EC: data = 12'h435;
        15'h02ED: data = 12'h439;
        15'h02EE: data = 12'h435;
        15'h02EF: data = 12'h433;
        15'h02F0: data = 12'h42F;
        15'h02F1: data = 12'h428;
        15'h02F2: data = 12'h42C;
        15'h02F3: data = 12'h42C;
        15'h02F4: data = 12'h42D;
        15'h02F5: data = 12'h432;
        15'h02F6: data = 12'h434;
        15'h02F7: data = 12'h438;
        15'h02F8: data = 12'h439;
        15'h02F9: data = 12'h432;
        15'h02FA: data = 12'h42B;
        15'h02FB: data = 12'h42A;
        15'h02FC: data = 12'h44A;
        15'h02FD: data = 12'h44C;
        15'h02FE: data = 12'h451;
        15'h02FF: data = 12'h456;
        15'h0300: data = 12'h456;
        15'h0301: data = 12'h456;
        15'h0302: data = 12'h455;
        15'h0303: data = 12'h44F;
        15'h0304: data = 12'h44B;
        15'h0305: data = 12'h447;
        15'h0306: data = 12'h44B;
        15'h0307: data = 12'h44D;
        15'h0308: data = 12'h453;
        15'h0309: data = 12'h455;
        15'h030A: data = 12'h453;
        15'h030B: data = 12'h451;
        15'h030C: data = 12'h44D;
        15'h030D: data = 12'h447;
        15'h030E: data = 12'h449;
        15'h030F: data = 12'h44C;
        15'h0310: data = 12'h44E;
        15'h0311: data = 12'h455;
        15'h0312: data = 12'h454;
        15'h0313: data = 12'h455;
        15'h0314: data = 12'h454;
        15'h0315: data = 12'h455;
        15'h0316: data = 12'h44C;
        15'h0317: data = 12'h44B;
        15'h0318: data = 12'h44C;
        15'h0319: data = 12'h44C;
        15'h031A: data = 12'h454;
        15'h031B: data = 12'h453;
        15'h031C: data = 12'h455;
        15'h031D: data = 12'h458;
        15'h031E: data = 12'h456;
        15'h031F: data = 12'h451;
        15'h0320: data = 12'h44B;
        15'h0321: data = 12'h44A;
        15'h0322: data = 12'h44B;
        15'h0323: data = 12'h450;
        15'h0324: data = 12'h452;
        15'h0325: data = 12'h455;
        15'h0326: data = 12'h454;
        15'h0327: data = 12'h454;
        15'h0328: data = 12'h44F;
        15'h0329: data = 12'h44B;
        15'h032A: data = 12'h447;
        15'h032B: data = 12'h44B;
        15'h032C: data = 12'h44F;
        15'h032D: data = 12'h456;
        15'h032E: data = 12'h457;
        15'h032F: data = 12'h455;
        15'h0330: data = 12'h457;
        15'h0331: data = 12'h452;
        15'h0332: data = 12'h44A;
        15'h0333: data = 12'h44C;
        15'h0334: data = 12'h44C;
        15'h0335: data = 12'h44F;
        15'h0336: data = 12'h455;
        15'h0337: data = 12'h456;
        15'h0338: data = 12'h456;
        15'h0339: data = 12'h457;
        15'h033A: data = 12'h450;
        15'h033B: data = 12'h44C;
        15'h033C: data = 12'h446;
        15'h033D: data = 12'h44A;
        15'h033E: data = 12'h449;
        15'h033F: data = 12'h456;
        15'h0340: data = 12'h456;
        15'h0341: data = 12'h456;
        15'h0342: data = 12'h453;
        15'h0343: data = 12'h451;
        15'h0344: data = 12'h44D;
        15'h0345: data = 12'h449;
        15'h0346: data = 12'h44B;
        15'h0347: data = 12'h44A;
        15'h0348: data = 12'h450;
        15'h0349: data = 12'h453;
        15'h034A: data = 12'h457;
        15'h034B: data = 12'h453;
        15'h034C: data = 12'h453;
        15'h034D: data = 12'h44D;
        15'h034E: data = 12'h44A;
        15'h034F: data = 12'h447;
        15'h0350: data = 12'h449;
        15'h0351: data = 12'h44C;
        15'h0352: data = 12'h452;
        15'h0353: data = 12'h456;
        15'h0354: data = 12'h457;
        15'h0355: data = 12'h457;
        15'h0356: data = 12'h455;
        15'h0357: data = 12'h44F;
        15'h0358: data = 12'h467;
        15'h0359: data = 12'h469;
        15'h035A: data = 12'h46A;
        15'h035B: data = 12'h46E;
        15'h035C: data = 12'h471;
        15'h035D: data = 12'h475;
        15'h035E: data = 12'h476;
        15'h035F: data = 12'h470;
        15'h0360: data = 12'h472;
        15'h0361: data = 12'h469;
        15'h0362: data = 12'h468;
        15'h0363: data = 12'h465;
        15'h0364: data = 12'h46B;
        15'h0365: data = 12'h46D;
        15'h0366: data = 12'h476;
        15'h0367: data = 12'h473;
        15'h0368: data = 12'h474;
        15'h0369: data = 12'h472;
        15'h036A: data = 12'h46B;
        15'h036B: data = 12'h469;
        15'h036C: data = 12'h465;
        15'h036D: data = 12'h468;
        15'h036E: data = 12'h46F;
        15'h036F: data = 12'h474;
        15'h0370: data = 12'h475;
        15'h0371: data = 12'h473;
        15'h0372: data = 12'h475;
        15'h0373: data = 12'h474;
        15'h0374: data = 12'h46B;
        15'h0375: data = 12'h46B;
        15'h0376: data = 12'h46E;
        15'h0377: data = 12'h46D;
        15'h0378: data = 12'h474;
        15'h0379: data = 12'h475;
        15'h037A: data = 12'h471;
        15'h037B: data = 12'h475;
        15'h037C: data = 12'h471;
        15'h037D: data = 12'h46D;
        15'h037E: data = 12'h46B;
        15'h037F: data = 12'h467;
        15'h0380: data = 12'h46B;
        15'h0381: data = 12'h470;
        15'h0382: data = 12'h472;
        15'h0383: data = 12'h473;
        15'h0384: data = 12'h477;
        15'h0385: data = 12'h471;
        15'h0386: data = 12'h473;
        15'h0387: data = 12'h46E;
        15'h0388: data = 12'h46A;
        15'h0389: data = 12'h468;
        15'h038A: data = 12'h46B;
        15'h038B: data = 12'h471;
        15'h038C: data = 12'h471;
        15'h038D: data = 12'h478;
        15'h038E: data = 12'h474;
        15'h038F: data = 12'h473;
        15'h0390: data = 12'h46D;
        15'h0391: data = 12'h46C;
        15'h0392: data = 12'h46B;
        15'h0393: data = 12'h46C;
        15'h0394: data = 12'h46F;
        15'h0395: data = 12'h471;
        15'h0396: data = 12'h473;
        15'h0397: data = 12'h473;
        15'h0398: data = 12'h475;
        15'h0399: data = 12'h46F;
        15'h039A: data = 12'h46B;
        15'h039B: data = 12'h46B;
        15'h039C: data = 12'h46C;
        15'h039D: data = 12'h46C;
        15'h039E: data = 12'h473;
        15'h039F: data = 12'h475;
        15'h03A0: data = 12'h472;
        15'h03A1: data = 12'h471;
        15'h03A2: data = 12'h470;
        15'h03A3: data = 12'h46D;
        15'h03A4: data = 12'h46A;
        15'h03A5: data = 12'h46B;
        15'h03A6: data = 12'h46B;
        15'h03A7: data = 12'h470;
        15'h03A8: data = 12'h474;
        15'h03A9: data = 12'h477;
        15'h03AA: data = 12'h477;
        15'h03AB: data = 12'h473;
        15'h03AC: data = 12'h46D;
        15'h03AD: data = 12'h469;
        15'h03AE: data = 12'h467;
        15'h03AF: data = 12'h468;
        15'h03B0: data = 12'h46A;
        15'h03B1: data = 12'h472;
        15'h03B2: data = 12'h473;
        15'h03B3: data = 12'h477;
        15'h03B4: data = 12'h49A;
        15'h03B5: data = 12'h48F;
        15'h03B6: data = 12'h48B;
        15'h03B7: data = 12'h487;
        15'h03B8: data = 12'h487;
        15'h03B9: data = 12'h488;
        15'h03BA: data = 12'h48E;
        15'h03BB: data = 12'h496;
        15'h03BC: data = 12'h499;
        15'h03BD: data = 12'h49B;
        15'h03BE: data = 12'h496;
        15'h03BF: data = 12'h48F;
        15'h03C0: data = 12'h489;
        15'h03C1: data = 12'h486;
        15'h03C2: data = 12'h489;
        15'h03C3: data = 12'h48F;
        15'h03C4: data = 12'h493;
        15'h03C5: data = 12'h498;
        15'h03C6: data = 12'h498;
        15'h03C7: data = 12'h496;
        15'h03C8: data = 12'h490;
        15'h03C9: data = 12'h48C;
        15'h03CA: data = 12'h486;
        15'h03CB: data = 12'h488;
        15'h03CC: data = 12'h48D;
        15'h03CD: data = 12'h48C;
        15'h03CE: data = 12'h494;
        15'h03CF: data = 12'h493;
        15'h03D0: data = 12'h497;
        15'h03D1: data = 12'h494;
        15'h03D2: data = 12'h48C;
        15'h03D3: data = 12'h487;
        15'h03D4: data = 12'h489;
        15'h03D5: data = 12'h489;
        15'h03D6: data = 12'h48D;
        15'h03D7: data = 12'h497;
        15'h03D8: data = 12'h495;
        15'h03D9: data = 12'h497;
        15'h03DA: data = 12'h494;
        15'h03DB: data = 12'h491;
        15'h03DC: data = 12'h48C;
        15'h03DD: data = 12'h48A;
        15'h03DE: data = 12'h48A;
        15'h03DF: data = 12'h490;
        15'h03E0: data = 12'h491;
        15'h03E1: data = 12'h498;
        15'h03E2: data = 12'h496;
        15'h03E3: data = 12'h49A;
        15'h03E4: data = 12'h493;
        15'h03E5: data = 12'h48C;
        15'h03E6: data = 12'h486;
        15'h03E7: data = 12'h487;
        15'h03E8: data = 12'h48D;
        15'h03E9: data = 12'h492;
        15'h03EA: data = 12'h494;
        15'h03EB: data = 12'h499;
        15'h03EC: data = 12'h493;
        15'h03ED: data = 12'h492;
        15'h03EE: data = 12'h490;
        15'h03EF: data = 12'h48E;
        15'h03F0: data = 12'h488;
        15'h03F1: data = 12'h48C;
        15'h03F2: data = 12'h48F;
        15'h03F3: data = 12'h493;
        15'h03F4: data = 12'h497;
        15'h03F5: data = 12'h495;
        15'h03F6: data = 12'h498;
        15'h03F7: data = 12'h492;
        15'h03F8: data = 12'h490;
        15'h03F9: data = 12'h48C;
        15'h03FA: data = 12'h48A;
        15'h03FB: data = 12'h48C;
        15'h03FC: data = 12'h491;
        15'h03FD: data = 12'h492;
        15'h03FE: data = 12'h496;
        15'h03FF: data = 12'h496;
        15'h0400: data = 12'h496;
        15'h0401: data = 12'h48F;
        15'h0402: data = 12'h491;
        15'h0403: data = 12'h4AC;
        15'h0404: data = 12'h4AB;
        15'h0405: data = 12'h4AF;
        15'h0406: data = 12'h4AC;
        15'h0407: data = 12'h4B3;
        15'h0408: data = 12'h4B4;
        15'h0409: data = 12'h4B5;
        15'h040A: data = 12'h4B6;
        15'h040B: data = 12'h4AB;
        15'h040C: data = 12'h4A9;
        15'h040D: data = 12'h4AC;
        15'h040E: data = 12'h4AD;
        15'h040F: data = 12'h4AB;
        15'h0410: data = 12'h4B4;
        15'h0411: data = 12'h4B5;
        15'h0412: data = 12'h4B5;
        15'h0413: data = 12'h4B6;
        15'h0414: data = 12'h4B1;
        15'h0415: data = 12'h4AE;
        15'h0416: data = 12'h4AD;
        15'h0417: data = 12'h4A7;
        15'h0418: data = 12'h4AD;
        15'h0419: data = 12'h4B1;
        15'h041A: data = 12'h4B9;
        15'h041B: data = 12'h4BC;
        15'h041C: data = 12'h4B8;
        15'h041D: data = 12'h4B4;
        15'h041E: data = 12'h4B1;
        15'h041F: data = 12'h4AE;
        15'h0420: data = 12'h4A8;
        15'h0421: data = 12'h4AB;
        15'h0422: data = 12'h4AE;
        15'h0423: data = 12'h4B6;
        15'h0424: data = 12'h4B9;
        15'h0425: data = 12'h4B8;
        15'h0426: data = 12'h4B3;
        15'h0427: data = 12'h4AF;
        15'h0428: data = 12'h4AA;
        15'h0429: data = 12'h4A5;
        15'h042A: data = 12'h4AB;
        15'h042B: data = 12'h4AD;
        15'h042C: data = 12'h4B0;
        15'h042D: data = 12'h4B6;
        15'h042E: data = 12'h4B7;
        15'h042F: data = 12'h4B7;
        15'h0430: data = 12'h4B1;
        15'h0431: data = 12'h4AC;
        15'h0432: data = 12'h4A8;
        15'h0433: data = 12'h4A8;
        15'h0434: data = 12'h4AB;
        15'h0435: data = 12'h4AE;
        15'h0436: data = 12'h4B6;
        15'h0437: data = 12'h4B5;
        15'h0438: data = 12'h4B5;
        15'h0439: data = 12'h4B6;
        15'h043A: data = 12'h4AD;
        15'h043B: data = 12'h4A8;
        15'h043C: data = 12'h4A8;
        15'h043D: data = 12'h4A7;
        15'h043E: data = 12'h4AB;
        15'h043F: data = 12'h4B4;
        15'h0440: data = 12'h4B3;
        15'h0441: data = 12'h4B4;
        15'h0442: data = 12'h4B0;
        15'h0443: data = 12'h4B0;
        15'h0444: data = 12'h4AC;
        15'h0445: data = 12'h4A9;
        15'h0446: data = 12'h4A9;
        15'h0447: data = 12'h4AA;
        15'h0448: data = 12'h4B1;
        15'h0449: data = 12'h4B5;
        15'h044A: data = 12'h4B5;
        15'h044B: data = 12'h4B5;
        15'h044C: data = 12'h4B3;
        15'h044D: data = 12'h4B0;
        15'h044E: data = 12'h4AD;
        15'h044F: data = 12'h4AB;
        15'h0450: data = 12'h4A7;
        15'h0451: data = 12'h4AC;
        15'h0452: data = 12'h4AF;
        15'h0453: data = 12'h4B6;
        15'h0454: data = 12'h4B9;
        15'h0455: data = 12'h4B5;
        15'h0456: data = 12'h4B3;
        15'h0457: data = 12'h4AD;
        15'h0458: data = 12'h4A6;
        15'h0459: data = 12'h4A5;
        15'h045A: data = 12'h4AA;
        15'h045B: data = 12'h4B0;
        15'h045C: data = 12'h4B8;
        15'h045D: data = 12'h4B9;
        15'h045E: data = 12'h4B7;
        15'h045F: data = 12'h4B5;
        15'h0460: data = 12'h4B3;
        15'h0461: data = 12'h4AA;
        15'h0462: data = 12'h4A4;
        15'h0463: data = 12'h4A9;
        15'h0464: data = 12'h4AC;
        15'h0465: data = 12'h4AE;
        15'h0466: data = 12'h4B5;
        15'h0467: data = 12'h4B5;
        15'h0468: data = 12'h4B5;
        15'h0469: data = 12'h4B5;
        15'h046A: data = 12'h4B0;
        15'h046B: data = 12'h4CA;
        15'h046C: data = 12'h4C6;
        15'h046D: data = 12'h4CE;
        15'h046E: data = 12'h4D0;
        15'h046F: data = 12'h4D3;
        15'h0470: data = 12'h4D8;
        15'h0471: data = 12'h4D4;
        15'h0472: data = 12'h4D5;
        15'h0473: data = 12'h4D4;
        15'h0474: data = 12'h4CD;
        15'h0475: data = 12'h4CB;
        15'h0476: data = 12'h4C9;
        15'h0477: data = 12'h4CC;
        15'h0478: data = 12'h4D1;
        15'h0479: data = 12'h4D5;
        15'h047A: data = 12'h4D6;
        15'h047B: data = 12'h4D8;
        15'h047C: data = 12'h4D1;
        15'h047D: data = 12'h4C9;
        15'h047E: data = 12'h4CA;
        15'h047F: data = 12'h4C9;
        15'h0480: data = 12'h4C6;
        15'h0481: data = 12'h4D1;
        15'h0482: data = 12'h4D3;
        15'h0483: data = 12'h4D5;
        15'h0484: data = 12'h4D5;
        15'h0485: data = 12'h4CF;
        15'h0486: data = 12'h4CD;
        15'h0487: data = 12'h4CA;
        15'h0488: data = 12'h4C9;
        15'h0489: data = 12'h4C9;
        15'h048A: data = 12'h4D0;
        15'h048B: data = 12'h4D1;
        15'h048C: data = 12'h4D7;
        15'h048D: data = 12'h4D7;
        15'h048E: data = 12'h4D5;
        15'h048F: data = 12'h4D3;
        15'h0490: data = 12'h4CB;
        15'h0491: data = 12'h4CA;
        15'h0492: data = 12'h4C7;
        15'h0493: data = 12'h4CF;
        15'h0494: data = 12'h4D0;
        15'h0495: data = 12'h4D5;
        15'h0496: data = 12'h4D8;
        15'h0497: data = 12'h4D4;
        15'h0498: data = 12'h4D8;
        15'h0499: data = 12'h4CF;
        15'h049A: data = 12'h4CC;
        15'h049B: data = 12'h4CA;
        15'h049C: data = 12'h4C9;
        15'h049D: data = 12'h4CE;
        15'h049E: data = 12'h4D4;
        15'h049F: data = 12'h4D9;
        15'h04A0: data = 12'h4D7;
        15'h04A1: data = 12'h4D5;
        15'h04A2: data = 12'h4CF;
        15'h04A3: data = 12'h4CC;
        15'h04A4: data = 12'h4CA;
        15'h04A5: data = 12'h4C9;
        15'h04A6: data = 12'h4C7;
        15'h04A7: data = 12'h4CE;
        15'h04A8: data = 12'h4D3;
        15'h04A9: data = 12'h4D9;
        15'h04AA: data = 12'h4D6;
        15'h04AB: data = 12'h4D5;
        15'h04AC: data = 12'h4CE;
        15'h04AD: data = 12'h4CE;
        15'h04AE: data = 12'h4C9;
        15'h04AF: data = 12'h4CD;
        15'h04B0: data = 12'h4CB;
        15'h04B1: data = 12'h4D0;
        15'h04B2: data = 12'h4D2;
        15'h04B3: data = 12'h4D5;
        15'h04B4: data = 12'h4D6;
        15'h04B5: data = 12'h4D2;
        15'h04B6: data = 12'h4CF;
        15'h04B7: data = 12'h4CD;
        15'h04B8: data = 12'h4CA;
        15'h04B9: data = 12'h4CE;
        15'h04BA: data = 12'h4CD;
        15'h04BB: data = 12'h4D6;
        15'h04BC: data = 12'h4D4;
        15'h04BD: data = 12'h4D8;
        15'h04BE: data = 12'h4D8;
        15'h04BF: data = 12'h4D2;
        15'h04C0: data = 12'h4CC;
        15'h04C1: data = 12'h4CD;
        15'h04C2: data = 12'h4CB;
        15'h04C3: data = 12'h4CB;
        15'h04C4: data = 12'h4D0;
        15'h04C5: data = 12'h4D3;
        15'h04C6: data = 12'h4D6;
        15'h04C7: data = 12'h4F4;
        15'h04C8: data = 12'h4F4;
        15'h04C9: data = 12'h4EF;
        15'h04CA: data = 12'h4E9;
        15'h04CB: data = 12'h4EA;
        15'h04CC: data = 12'h4EC;
        15'h04CD: data = 12'h4EF;
        15'h04CE: data = 12'h4F4;
        15'h04CF: data = 12'h4F6;
        15'h04D0: data = 12'h4F5;
        15'h04D1: data = 12'h4F5;
        15'h04D2: data = 12'h4EE;
        15'h04D3: data = 12'h4EA;
        15'h04D4: data = 12'h4E9;
        15'h04D5: data = 12'h4E9;
        15'h04D6: data = 12'h4EC;
        15'h04D7: data = 12'h4F2;
        15'h04D8: data = 12'h4F9;
        15'h04D9: data = 12'h4F6;
        15'h04DA: data = 12'h4FA;
        15'h04DB: data = 12'h4F2;
        15'h04DC: data = 12'h4EC;
        15'h04DD: data = 12'h4EB;
        15'h04DE: data = 12'h4EB;
        15'h04DF: data = 12'h4EA;
        15'h04E0: data = 12'h4F3;
        15'h04E1: data = 12'h4F6;
        15'h04E2: data = 12'h4FB;
        15'h04E3: data = 12'h4F6;
        15'h04E4: data = 12'h4F6;
        15'h04E5: data = 12'h4F2;
        15'h04E6: data = 12'h4EC;
        15'h04E7: data = 12'h4E9;
        15'h04E8: data = 12'h4EC;
        15'h04E9: data = 12'h4F1;
        15'h04EA: data = 12'h4F6;
        15'h04EB: data = 12'h4F7;
        15'h04EC: data = 12'h4F6;
        15'h04ED: data = 12'h4F7;
        15'h04EE: data = 12'h4F3;
        15'h04EF: data = 12'h4EE;
        15'h04F0: data = 12'h4EE;
        15'h04F1: data = 12'h4ED;
        15'h04F2: data = 12'h4F0;
        15'h04F3: data = 12'h4F3;
        15'h04F4: data = 12'h4F9;
        15'h04F5: data = 12'h4F8;
        15'h04F6: data = 12'h4F5;
        15'h04F7: data = 12'h4F7;
        15'h04F8: data = 12'h4F2;
        15'h04F9: data = 12'h4ED;
        15'h04FA: data = 12'h4E7;
        15'h04FB: data = 12'h4EA;
        15'h04FC: data = 12'h4EC;
        15'h04FD: data = 12'h4F3;
        15'h04FE: data = 12'h4F4;
        15'h04FF: data = 12'h4F9;
        15'h0500: data = 12'h4F8;
        15'h0501: data = 12'h4F5;
        15'h0502: data = 12'h4F0;
        15'h0503: data = 12'h4EA;
        15'h0504: data = 12'h4E9;
        15'h0505: data = 12'h4EC;
        15'h0506: data = 12'h4F0;
        15'h0507: data = 12'h4F3;
        15'h0508: data = 12'h4F7;
        15'h0509: data = 12'h4F5;
        15'h050A: data = 12'h4F5;
        15'h050B: data = 12'h4F1;
        15'h050C: data = 12'h4EC;
        15'h050D: data = 12'h4E6;
        15'h050E: data = 12'h4EA;
        15'h050F: data = 12'h4EC;
        15'h0510: data = 12'h4F3;
        15'h0511: data = 12'h4F5;
        15'h0512: data = 12'h4F9;
        15'h0513: data = 12'h4F7;
        15'h0514: data = 12'h4F2;
        15'h0515: data = 12'h4EC;
        15'h0516: data = 12'h50A;
        15'h0517: data = 12'h50C;
        15'h0518: data = 12'h50F;
        15'h0519: data = 12'h50E;
        15'h051A: data = 12'h515;
        15'h051B: data = 12'h515;
        15'h051C: data = 12'h513;
        15'h051D: data = 12'h514;
        15'h051E: data = 12'h50E;
        15'h051F: data = 12'h50F;
        15'h0520: data = 12'h50A;
        15'h0521: data = 12'h50A;
        15'h0522: data = 12'h50E;
        15'h0523: data = 12'h512;
        15'h0524: data = 12'h515;
        15'h0525: data = 12'h51A;
        15'h0526: data = 12'h517;
        15'h0527: data = 12'h517;
        15'h0528: data = 12'h50F;
        15'h0529: data = 12'h50C;
        15'h052A: data = 12'h50B;
        15'h052B: data = 12'h511;
        15'h052C: data = 12'h512;
        15'h052D: data = 12'h513;
        15'h052E: data = 12'h517;
        15'h052F: data = 12'h51D;
        15'h0530: data = 12'h518;
        15'h0531: data = 12'h516;
        15'h0532: data = 12'h50F;
        15'h0533: data = 12'h50F;
        15'h0534: data = 12'h50D;
        15'h0535: data = 12'h512;
        15'h0536: data = 12'h517;
        15'h0537: data = 12'h515;
        15'h0538: data = 12'h517;
        15'h0539: data = 12'h514;
        15'h053A: data = 12'h513;
        15'h053B: data = 12'h50F;
        15'h053C: data = 12'h50D;
        15'h053D: data = 12'h50C;
        15'h053E: data = 12'h50E;
        15'h053F: data = 12'h510;
        15'h0540: data = 12'h514;
        15'h0541: data = 12'h517;
        15'h0542: data = 12'h519;
        15'h0543: data = 12'h517;
        15'h0544: data = 12'h513;
        15'h0545: data = 12'h50F;
        15'h0546: data = 12'h50D;
        15'h0547: data = 12'h50E;
        15'h0548: data = 12'h50F;
        15'h0549: data = 12'h515;
        15'h054A: data = 12'h51A;
        15'h054B: data = 12'h51B;
        15'h054C: data = 12'h517;
        15'h054D: data = 12'h516;
        15'h054E: data = 12'h50F;
        15'h054F: data = 12'h50E;
        15'h0550: data = 12'h50E;
        15'h0551: data = 12'h50D;
        15'h0552: data = 12'h511;
        15'h0553: data = 12'h512;
        15'h0554: data = 12'h514;
        15'h0555: data = 12'h516;
        15'h0556: data = 12'h517;
        15'h0557: data = 12'h514;
        15'h0558: data = 12'h50B;
        15'h0559: data = 12'h50D;
        15'h055A: data = 12'h50A;
        15'h055B: data = 12'h50F;
        15'h055C: data = 12'h512;
        15'h055D: data = 12'h518;
        15'h055E: data = 12'h515;
        15'h055F: data = 12'h515;
        15'h0560: data = 12'h516;
        15'h0561: data = 12'h511;
        15'h0562: data = 12'h50D;
        15'h0563: data = 12'h50B;
        15'h0564: data = 12'h50A;
        15'h0565: data = 12'h50E;
        15'h0566: data = 12'h513;
        15'h0567: data = 12'h515;
        15'h0568: data = 12'h511;
        15'h0569: data = 12'h517;
        15'h056A: data = 12'h510;
        15'h056B: data = 12'h50D;
        15'h056C: data = 12'h50D;
        15'h056D: data = 12'h509;
        15'h056E: data = 12'h50C;
        15'h056F: data = 12'h513;
        15'h0570: data = 12'h513;
        15'h0571: data = 12'h522;
        15'h0572: data = 12'h52D;
        15'h0573: data = 12'h526;
        15'h0574: data = 12'h522;
        15'h0575: data = 12'h523;
        15'h0576: data = 12'h51C;
        15'h0577: data = 12'h522;
        15'h0578: data = 12'h524;
        15'h0579: data = 12'h52B;
        15'h057A: data = 12'h52D;
        15'h057B: data = 12'h52D;
        15'h057C: data = 12'h52B;
        15'h057D: data = 12'h527;
        15'h057E: data = 12'h51E;
        15'h057F: data = 12'h51D;
        15'h0580: data = 12'h521;
        15'h0581: data = 12'h524;
        15'h0582: data = 12'h52B;
        15'h0583: data = 12'h52D;
        15'h0584: data = 12'h52D;
        15'h0585: data = 12'h52E;
        15'h0586: data = 12'h524;
        15'h0587: data = 12'h51E;
        15'h0588: data = 12'h51F;
        15'h0589: data = 12'h51C;
        15'h058A: data = 12'h522;
        15'h058B: data = 12'h52A;
        15'h058C: data = 12'h52B;
        15'h058D: data = 12'h52F;
        15'h058E: data = 12'h52B;
        15'h058F: data = 12'h525;
        15'h0590: data = 12'h51E;
        15'h0591: data = 12'h51C;
        15'h0592: data = 12'h51D;
        15'h0593: data = 12'h522;
        15'h0594: data = 12'h524;
        15'h0595: data = 12'h52A;
        15'h0596: data = 12'h52C;
        15'h0597: data = 12'h52B;
        15'h0598: data = 12'h529;
        15'h0599: data = 12'h526;
        15'h059A: data = 12'h51E;
        15'h059B: data = 12'h51E;
        15'h059C: data = 12'h51E;
        15'h059D: data = 12'h520;
        15'h059E: data = 12'h529;
        15'h059F: data = 12'h52C;
        15'h05A0: data = 12'h52D;
        15'h05A1: data = 12'h52D;
        15'h05A2: data = 12'h528;
        15'h05A3: data = 12'h51E;
        15'h05A4: data = 12'h51C;
        15'h05A5: data = 12'h51C;
        15'h05A6: data = 12'h523;
        15'h05A7: data = 12'h524;
        15'h05A8: data = 12'h529;
        15'h05A9: data = 12'h528;
        15'h05AA: data = 12'h527;
        15'h05AB: data = 12'h526;
        15'h05AC: data = 12'h520;
        15'h05AD: data = 12'h51B;
        15'h05AE: data = 12'h520;
        15'h05AF: data = 12'h521;
        15'h05B0: data = 12'h523;
        15'h05B1: data = 12'h529;
        15'h05B2: data = 12'h52E;
        15'h05B3: data = 12'h52A;
        15'h05B4: data = 12'h52A;
        15'h05B5: data = 12'h522;
        15'h05B6: data = 12'h51F;
        15'h05B7: data = 12'h520;
        15'h05B8: data = 12'h521;
        15'h05B9: data = 12'h525;
        15'h05BA: data = 12'h528;
        15'h05BB: data = 12'h52A;
        15'h05BC: data = 12'h528;
        15'h05BD: data = 12'h529;
        15'h05BE: data = 12'h523;
        15'h05BF: data = 12'h520;
        15'h05C0: data = 12'h542;
        15'h05C1: data = 12'h541;
        15'h05C2: data = 12'h542;
        15'h05C3: data = 12'h547;
        15'h05C4: data = 12'h546;
        15'h05C5: data = 12'h549;
        15'h05C6: data = 12'h545;
        15'h05C7: data = 12'h546;
        15'h05C8: data = 12'h543;
        15'h05C9: data = 12'h542;
        15'h05CA: data = 12'h53C;
        15'h05CB: data = 12'h540;
        15'h05CC: data = 12'h541;
        15'h05CD: data = 12'h547;
        15'h05CE: data = 12'h54C;
        15'h05CF: data = 12'h54D;
        15'h05D0: data = 12'h54C;
        15'h05D1: data = 12'h548;
        15'h05D2: data = 12'h542;
        15'h05D3: data = 12'h53A;
        15'h05D4: data = 12'h540;
        15'h05D5: data = 12'h542;
        15'h05D6: data = 12'h548;
        15'h05D7: data = 12'h54B;
        15'h05D8: data = 12'h54C;
        15'h05D9: data = 12'h548;
        15'h05DA: data = 12'h549;
        15'h05DB: data = 12'h541;
        15'h05DC: data = 12'h53C;
        15'h05DD: data = 12'h53E;
        15'h05DE: data = 12'h542;
        15'h05DF: data = 12'h543;
        15'h05E0: data = 12'h54B;
        15'h05E1: data = 12'h54C;
        15'h05E2: data = 12'h54A;
        15'h05E3: data = 12'h54B;
        15'h05E4: data = 12'h544;
        15'h05E5: data = 12'h53F;
        15'h05E6: data = 12'h53E;
        15'h05E7: data = 12'h542;
        15'h05E8: data = 12'h543;
        15'h05E9: data = 12'h549;
        15'h05EA: data = 12'h54B;
        15'h05EB: data = 12'h54D;
        15'h05EC: data = 12'h54B;
        15'h05ED: data = 12'h545;
        15'h05EE: data = 12'h53F;
        15'h05EF: data = 12'h53F;
        15'h05F0: data = 12'h53B;
        15'h05F1: data = 12'h541;
        15'h05F2: data = 12'h545;
        15'h05F3: data = 12'h549;
        15'h05F4: data = 12'h549;
        15'h05F5: data = 12'h549;
        15'h05F6: data = 12'h546;
        15'h05F7: data = 12'h543;
        15'h05F8: data = 12'h53D;
        15'h05F9: data = 12'h540;
        15'h05FA: data = 12'h541;
        15'h05FB: data = 12'h544;
        15'h05FC: data = 12'h54A;
        15'h05FD: data = 12'h549;
        15'h05FE: data = 12'h54A;
        15'h05FF: data = 12'h547;
        15'h0600: data = 12'h547;
        15'h0601: data = 12'h542;
        15'h0602: data = 12'h53E;
        15'h0603: data = 12'h53E;
        15'h0604: data = 12'h53D;
        15'h0605: data = 12'h544;
        15'h0606: data = 12'h547;
        15'h0607: data = 12'h548;
        15'h0608: data = 12'h546;
        15'h0609: data = 12'h546;
        15'h060A: data = 12'h545;
        15'h060B: data = 12'h542;
        15'h060C: data = 12'h53C;
        15'h060D: data = 12'h541;
        15'h060E: data = 12'h547;
        15'h060F: data = 12'h56C;
        15'h0610: data = 12'h568;
        15'h0611: data = 12'h569;
        15'h0612: data = 12'h56A;
        15'h0613: data = 12'h566;
        15'h0614: data = 12'h563;
        15'h0615: data = 12'h55F;
        15'h0616: data = 12'h561;
        15'h0617: data = 12'h562;
        15'h0618: data = 12'h564;
        15'h0619: data = 12'h568;
        15'h061A: data = 12'h56A;
        15'h061B: data = 12'h56C;
        15'h061C: data = 12'h568;
        15'h061D: data = 12'h567;
        15'h061E: data = 12'h55F;
        15'h061F: data = 12'h55F;
        15'h0620: data = 12'h560;
        15'h0621: data = 12'h562;
        15'h0622: data = 12'h569;
        15'h0623: data = 12'h56E;
        15'h0624: data = 12'h56D;
        15'h0625: data = 12'h568;
        15'h0626: data = 12'h566;
        15'h0627: data = 12'h564;
        15'h0628: data = 12'h560;
        15'h0629: data = 12'h55F;
        15'h062A: data = 12'h562;
        15'h062B: data = 12'h568;
        15'h062C: data = 12'h56B;
        15'h062D: data = 12'h56C;
        15'h062E: data = 12'h56A;
        15'h062F: data = 12'h569;
        15'h0630: data = 12'h565;
        15'h0631: data = 12'h560;
        15'h0632: data = 12'h55E;
        15'h0633: data = 12'h55F;
        15'h0634: data = 12'h566;
        15'h0635: data = 12'h569;
        15'h0636: data = 12'h56C;
        15'h0637: data = 12'h56F;
        15'h0638: data = 12'h569;
        15'h0639: data = 12'h565;
        15'h063A: data = 12'h562;
        15'h063B: data = 12'h561;
        15'h063C: data = 12'h561;
        15'h063D: data = 12'h564;
        15'h063E: data = 12'h56A;
        15'h063F: data = 12'h56A;
        15'h0640: data = 12'h569;
        15'h0641: data = 12'h567;
        15'h0642: data = 12'h56A;
        15'h0643: data = 12'h56A;
        15'h0644: data = 12'h562;
        15'h0645: data = 12'h563;
        15'h0646: data = 12'h561;
        15'h0647: data = 12'h566;
        15'h0648: data = 12'h56B;
        15'h0649: data = 12'h569;
        15'h064A: data = 12'h568;
        15'h064B: data = 12'h569;
        15'h064C: data = 12'h569;
        15'h064D: data = 12'h560;
        15'h064E: data = 12'h560;
        15'h064F: data = 12'h563;
        15'h0650: data = 12'h562;
        15'h0651: data = 12'h566;
        15'h0652: data = 12'h56B;
        15'h0653: data = 12'h571;
        15'h0654: data = 12'h56A;
        15'h0655: data = 12'h56B;
        15'h0656: data = 12'h564;
        15'h0657: data = 12'h561;
        15'h0658: data = 12'h562;
        15'h0659: data = 12'h562;
        15'h065A: data = 12'h569;
        15'h065B: data = 12'h570;
        15'h065C: data = 12'h56C;
        15'h065D: data = 12'h56B;
        15'h065E: data = 12'h569;
        15'h065F: data = 12'h562;
        15'h0660: data = 12'h561;
        15'h0661: data = 12'h560;
        15'h0662: data = 12'h564;
        15'h0663: data = 12'h566;
        15'h0664: data = 12'h569;
        15'h0665: data = 12'h56C;
        15'h0666: data = 12'h56C;
        15'h0667: data = 12'h569;
        15'h0668: data = 12'h567;
        15'h0669: data = 12'h564;
        15'h066A: data = 12'h565;
        15'h066B: data = 12'h563;
        15'h066C: data = 12'h565;
        15'h066D: data = 12'h56B;
        15'h066E: data = 12'h56A;
        15'h066F: data = 12'h56C;
        15'h0670: data = 12'h56B;
        15'h0671: data = 12'h569;
        15'h0672: data = 12'h566;
        15'h0673: data = 12'h563;
        15'h0674: data = 12'h562;
        15'h0675: data = 12'h562;
        15'h0676: data = 12'h567;
        15'h0677: data = 12'h56B;
        15'h0678: data = 12'h58E;
        15'h0679: data = 12'h58A;
        15'h067A: data = 12'h58B;
        15'h067B: data = 12'h586;
        15'h067C: data = 12'h582;
        15'h067D: data = 12'h57F;
        15'h067E: data = 12'h580;
        15'h067F: data = 12'h582;
        15'h0680: data = 12'h586;
        15'h0681: data = 12'h589;
        15'h0682: data = 12'h58C;
        15'h0683: data = 12'h58C;
        15'h0684: data = 12'h58A;
        15'h0685: data = 12'h586;
        15'h0686: data = 12'h580;
        15'h0687: data = 12'h57D;
        15'h0688: data = 12'h57F;
        15'h0689: data = 12'h57F;
        15'h068A: data = 12'h589;
        15'h068B: data = 12'h58F;
        15'h068C: data = 12'h58D;
        15'h068D: data = 12'h586;
        15'h068E: data = 12'h587;
        15'h068F: data = 12'h57D;
        15'h0690: data = 12'h57F;
        15'h0691: data = 12'h57D;
        15'h0692: data = 12'h581;
        15'h0693: data = 12'h58B;
        15'h0694: data = 12'h58A;
        15'h0695: data = 12'h58B;
        15'h0696: data = 12'h588;
        15'h0697: data = 12'h585;
        15'h0698: data = 12'h585;
        15'h0699: data = 12'h57F;
        15'h069A: data = 12'h57F;
        15'h069B: data = 12'h583;
        15'h069C: data = 12'h585;
        15'h069D: data = 12'h588;
        15'h069E: data = 12'h58B;
        15'h069F: data = 12'h58B;
        15'h06A0: data = 12'h588;
        15'h06A1: data = 12'h584;
        15'h06A2: data = 12'h580;
        15'h06A3: data = 12'h57C;
        15'h06A4: data = 12'h583;
        15'h06A5: data = 12'h582;
        15'h06A6: data = 12'h586;
        15'h06A7: data = 12'h586;
        15'h06A8: data = 12'h58C;
        15'h06A9: data = 12'h588;
        15'h06AA: data = 12'h588;
        15'h06AB: data = 12'h583;
        15'h06AC: data = 12'h57F;
        15'h06AD: data = 12'h580;
        15'h06AE: data = 12'h582;
        15'h06AF: data = 12'h583;
        15'h06B0: data = 12'h588;
        15'h06B1: data = 12'h589;
        15'h06B2: data = 12'h589;
        15'h06B3: data = 12'h58A;
        15'h06B4: data = 12'h586;
        15'h06B5: data = 12'h582;
        15'h06B6: data = 12'h57F;
        15'h06B7: data = 12'h57E;
        15'h06B8: data = 12'h581;
        15'h06B9: data = 12'h585;
        15'h06BA: data = 12'h588;
        15'h06BB: data = 12'h58A;
        15'h06BC: data = 12'h589;
        15'h06BD: data = 12'h586;
        15'h06BE: data = 12'h582;
        15'h06BF: data = 12'h585;
        15'h06C0: data = 12'h57D;
        15'h06C1: data = 12'h582;
        15'h06C2: data = 12'h585;
        15'h06C3: data = 12'h588;
        15'h06C4: data = 12'h58B;
        15'h06C5: data = 12'h58B;
        15'h06C6: data = 12'h5AC;
        15'h06C7: data = 12'h5AA;
        15'h06C8: data = 12'h5A3;
        15'h06C9: data = 12'h59F;
        15'h06CA: data = 12'h59B;
        15'h06CB: data = 12'h59F;
        15'h06CC: data = 12'h5A7;
        15'h06CD: data = 12'h5A8;
        15'h06CE: data = 12'h5AB;
        15'h06CF: data = 12'h5AB;
        15'h06D0: data = 12'h5A8;
        15'h06D1: data = 12'h5A6;
        15'h06D2: data = 12'h5A1;
        15'h06D3: data = 12'h59C;
        15'h06D4: data = 12'h59E;
        15'h06D5: data = 12'h59F;
        15'h06D6: data = 12'h5A7;
        15'h06D7: data = 12'h5AB;
        15'h06D8: data = 12'h5AA;
        15'h06D9: data = 12'h5AC;
        15'h06DA: data = 12'h5AA;
        15'h06DB: data = 12'h5A2;
        15'h06DC: data = 12'h59D;
        15'h06DD: data = 12'h5A1;
        15'h06DE: data = 12'h5A1;
        15'h06DF: data = 12'h5A5;
        15'h06E0: data = 12'h5A3;
        15'h06E1: data = 12'h5A9;
        15'h06E2: data = 12'h5AD;
        15'h06E3: data = 12'h5A9;
        15'h06E4: data = 12'h5A6;
        15'h06E5: data = 12'h59E;
        15'h06E6: data = 12'h59E;
        15'h06E7: data = 12'h59D;
        15'h06E8: data = 12'h5A0;
        15'h06E9: data = 12'h5A5;
        15'h06EA: data = 12'h5AE;
        15'h06EB: data = 12'h5AA;
        15'h06EC: data = 12'h5A7;
        15'h06ED: data = 12'h5A6;
        15'h06EE: data = 12'h59E;
        15'h06EF: data = 12'h59E;
        15'h06F0: data = 12'h59D;
        15'h06F1: data = 12'h59F;
        15'h06F2: data = 12'h5A5;
        15'h06F3: data = 12'h5AB;
        15'h06F4: data = 12'h5AD;
        15'h06F5: data = 12'h5AA;
        15'h06F6: data = 12'h5AA;
        15'h06F7: data = 12'h5A5;
        15'h06F8: data = 12'h5A2;
        15'h06F9: data = 12'h59B;
        15'h06FA: data = 12'h59F;
        15'h06FB: data = 12'h5A0;
        15'h06FC: data = 12'h5A8;
        15'h06FD: data = 12'h5A7;
        15'h06FE: data = 12'h5AC;
        15'h06FF: data = 12'h5A8;
        15'h0700: data = 12'h5A6;
        15'h0701: data = 12'h5A0;
        15'h0702: data = 12'h59E;
        15'h0703: data = 12'h5A0;
        15'h0704: data = 12'h5A1;
        15'h0705: data = 12'h5A6;
        15'h0706: data = 12'h5AD;
        15'h0707: data = 12'h5AD;
        15'h0708: data = 12'h5A9;
        15'h0709: data = 12'h5A6;
        15'h070A: data = 12'h5A1;
        15'h070B: data = 12'h59C;
        15'h070C: data = 12'h59F;
        15'h070D: data = 12'h59F;
        15'h070E: data = 12'h5A0;
        15'h070F: data = 12'h5A6;
        15'h0710: data = 12'h5AA;
        15'h0711: data = 12'h5A9;
        15'h0712: data = 12'h5AC;
        15'h0713: data = 12'h5A5;
        15'h0714: data = 12'h5A0;
        15'h0715: data = 12'h5C0;
        15'h0716: data = 12'h5BF;
        15'h0717: data = 12'h5C2;
        15'h0718: data = 12'h5C9;
        15'h0719: data = 12'h5CB;
        15'h071A: data = 12'h5CF;
        15'h071B: data = 12'h5C8;
        15'h071C: data = 12'h5C7;
        15'h071D: data = 12'h5C4;
        15'h071E: data = 12'h5BF;
        15'h071F: data = 12'h5C0;
        15'h0720: data = 12'h5BE;
        15'h0721: data = 12'h5C7;
        15'h0722: data = 12'h5CB;
        15'h0723: data = 12'h5CD;
        15'h0724: data = 12'h5CC;
        15'h0725: data = 12'h5CB;
        15'h0726: data = 12'h5C4;
        15'h0727: data = 12'h5BC;
        15'h0728: data = 12'h5BC;
        15'h0729: data = 12'h5BB;
        15'h072A: data = 12'h5C6;
        15'h072B: data = 12'h5CB;
        15'h072C: data = 12'h5CB;
        15'h072D: data = 12'h5CC;
        15'h072E: data = 12'h5CD;
        15'h072F: data = 12'h5C7;
        15'h0730: data = 12'h5C0;
        15'h0731: data = 12'h5BF;
        15'h0732: data = 12'h5C0;
        15'h0733: data = 12'h5BF;
        15'h0734: data = 12'h5C1;
        15'h0735: data = 12'h5C8;
        15'h0736: data = 12'h5C9;
        15'h0737: data = 12'h5CB;
        15'h0738: data = 12'h5CA;
        15'h0739: data = 12'h5C2;
        15'h073A: data = 12'h5C1;
        15'h073B: data = 12'h5C0;
        15'h073C: data = 12'h5BC;
        15'h073D: data = 12'h5C6;
        15'h073E: data = 12'h5C5;
        15'h073F: data = 12'h5CA;
        15'h0740: data = 12'h5C9;
        15'h0741: data = 12'h5C9;
        15'h0742: data = 12'h5C8;
        15'h0743: data = 12'h5C1;
        15'h0744: data = 12'h5C0;
        15'h0745: data = 12'h5BC;
        15'h0746: data = 12'h5BF;
        15'h0747: data = 12'h5C3;
        15'h0748: data = 12'h5C9;
        15'h0749: data = 12'h5CB;
        15'h074A: data = 12'h5CC;
        15'h074B: data = 12'h5CF;
        15'h074C: data = 12'h5C9;
        15'h074D: data = 12'h5C3;
        15'h074E: data = 12'h5BD;
        15'h074F: data = 12'h5BF;
        15'h0750: data = 12'h5C0;
        15'h0751: data = 12'h5C2;
        15'h0752: data = 12'h5CC;
        15'h0753: data = 12'h5C7;
        15'h0754: data = 12'h5CA;
        15'h0755: data = 12'h5C6;
        15'h0756: data = 12'h5C3;
        15'h0757: data = 12'h5BD;
        15'h0758: data = 12'h5BC;
        15'h0759: data = 12'h5BF;
        15'h075A: data = 12'h5C1;
        15'h075B: data = 12'h5C9;
        15'h075C: data = 12'h5CB;
        15'h075D: data = 12'h5CD;
        15'h075E: data = 12'h5CC;
        15'h075F: data = 12'h5CA;
        15'h0760: data = 12'h5C7;
        15'h0761: data = 12'h5C3;
        15'h0762: data = 12'h5BF;
        15'h0763: data = 12'h5C8;
        15'h0764: data = 12'h5E1;
        15'h0765: data = 12'h5EA;
        15'h0766: data = 12'h5EB;
        15'h0767: data = 12'h5EB;
        15'h0768: data = 12'h5ED;
        15'h0769: data = 12'h5E6;
        15'h076A: data = 12'h5E2;
        15'h076B: data = 12'h5DF;
        15'h076C: data = 12'h5E0;
        15'h076D: data = 12'h5E3;
        15'h076E: data = 12'h5E0;
        15'h076F: data = 12'h5E5;
        15'h0770: data = 12'h5EC;
        15'h0771: data = 12'h5E9;
        15'h0772: data = 12'h5E5;
        15'h0773: data = 12'h5E3;
        15'h0774: data = 12'h5E3;
        15'h0775: data = 12'h5E2;
        15'h0776: data = 12'h5E4;
        15'h0777: data = 12'h5E8;
        15'h0778: data = 12'h5EC;
        15'h0779: data = 12'h5EE;
        15'h077A: data = 12'h5EE;
        15'h077B: data = 12'h5ED;
        15'h077C: data = 12'h5E3;
        15'h077D: data = 12'h5E0;
        15'h077E: data = 12'h5DA;
        15'h077F: data = 12'h5DE;
        15'h0780: data = 12'h5E2;
        15'h0781: data = 12'h5E4;
        15'h0782: data = 12'h5EC;
        15'h0783: data = 12'h5EB;
        15'h0784: data = 12'h5EC;
        15'h0785: data = 12'h5E9;
        15'h0786: data = 12'h5E5;
        15'h0787: data = 12'h5E1;
        15'h0788: data = 12'h5E1;
        15'h0789: data = 12'h5E0;
        15'h078A: data = 12'h5E8;
        15'h078B: data = 12'h5EB;
        15'h078C: data = 12'h5ED;
        15'h078D: data = 12'h5EB;
        15'h078E: data = 12'h5EB;
        15'h078F: data = 12'h5E3;
        15'h0790: data = 12'h5E0;
        15'h0791: data = 12'h5E0;
        15'h0792: data = 12'h5E3;
        15'h0793: data = 12'h5E8;
        15'h0794: data = 12'h5EC;
        15'h0795: data = 12'h5F0;
        15'h0796: data = 12'h5EC;
        15'h0797: data = 12'h5EB;
        15'h0798: data = 12'h5E8;
        15'h0799: data = 12'h5E0;
        15'h079A: data = 12'h5DE;
        15'h079B: data = 12'h5DE;
        15'h079C: data = 12'h5E1;
        15'h079D: data = 12'h5E6;
        15'h079E: data = 12'h5E6;
        15'h079F: data = 12'h5EB;
        15'h07A0: data = 12'h5E7;
        15'h07A1: data = 12'h5E9;
        15'h07A2: data = 12'h5E6;
        15'h07A3: data = 12'h5E2;
        15'h07A4: data = 12'h5DF;
        15'h07A5: data = 12'h5E1;
        15'h07A6: data = 12'h5E4;
        15'h07A7: data = 12'h5EC;
        15'h07A8: data = 12'h5EE;
        15'h07A9: data = 12'h5EA;
        15'h07AA: data = 12'h5EB;
        15'h07AB: data = 12'h5E6;
        15'h07AC: data = 12'h5E3;
        15'h07AD: data = 12'h5E1;
        15'h07AE: data = 12'h5E1;
        15'h07AF: data = 12'h5E3;
        15'h07B0: data = 12'h5E6;
        15'h07B1: data = 12'h5EC;
        15'h07B2: data = 12'h60B;
        15'h07B3: data = 12'h610;
        15'h07B4: data = 12'h609;
        15'h07B5: data = 12'h608;
        15'h07B6: data = 12'h600;
        15'h07B7: data = 12'h5FF;
        15'h07B8: data = 12'h601;
        15'h07B9: data = 12'h603;
        15'h07BA: data = 12'h608;
        15'h07BB: data = 12'h60B;
        15'h07BC: data = 12'h60A;
        15'h07BD: data = 12'h60B;
        15'h07BE: data = 12'h608;
        15'h07BF: data = 12'h606;
        15'h07C0: data = 12'h5FF;
        15'h07C1: data = 12'h601;
        15'h07C2: data = 12'h5FF;
        15'h07C3: data = 12'h604;
        15'h07C4: data = 12'h605;
        15'h07C5: data = 12'h60D;
        15'h07C6: data = 12'h611;
        15'h07C7: data = 12'h60C;
        15'h07C8: data = 12'h609;
        15'h07C9: data = 12'h605;
        15'h07CA: data = 12'h603;
        15'h07CB: data = 12'h603;
        15'h07CC: data = 12'h603;
        15'h07CD: data = 12'h605;
        15'h07CE: data = 12'h60C;
        15'h07CF: data = 12'h60A;
        15'h07D0: data = 12'h60B;
        15'h07D1: data = 12'h60C;
        15'h07D2: data = 12'h606;
        15'h07D3: data = 12'h600;
        15'h07D4: data = 12'h600;
        15'h07D5: data = 12'h602;
        15'h07D6: data = 12'h605;
        15'h07D7: data = 12'h60D;
        15'h07D8: data = 12'h60B;
        15'h07D9: data = 12'h60F;
        15'h07DA: data = 12'h60D;
        15'h07DB: data = 12'h606;
        15'h07DC: data = 12'h605;
        15'h07DD: data = 12'h600;
        15'h07DE: data = 12'h5FD;
        15'h07DF: data = 12'h5FE;
        15'h07E0: data = 12'h603;
        15'h07E1: data = 12'h607;
        15'h07E2: data = 12'h60C;
        15'h07E3: data = 12'h60C;
        15'h07E4: data = 12'h60E;
        15'h07E5: data = 12'h609;
        15'h07E6: data = 12'h601;
        15'h07E7: data = 12'h5FE;
        15'h07E8: data = 12'h5FE;
        15'h07E9: data = 12'h5FF;
        15'h07EA: data = 12'h606;
        15'h07EB: data = 12'h60B;
        15'h07EC: data = 12'h60C;
        15'h07ED: data = 12'h60E;
        15'h07EE: data = 12'h60B;
        15'h07EF: data = 12'h603;
        15'h07F0: data = 12'h602;
        15'h07F1: data = 12'h601;
        15'h07F2: data = 12'h605;
        15'h07F3: data = 12'h600;
        15'h07F4: data = 12'h60C;
        15'h07F5: data = 12'h60C;
        15'h07F6: data = 12'h609;
        15'h07F7: data = 12'h609;
        15'h07F8: data = 12'h606;
        15'h07F9: data = 12'h603;
        15'h07FA: data = 12'h5FF;
        15'h07FB: data = 12'h5FF;
        15'h07FC: data = 12'h603;
        15'h07FD: data = 12'h607;
        15'h07FE: data = 12'h60C;
        15'h07FF: data = 12'h60B;
        15'h0800: data = 12'h607;
        15'h0801: data = 12'h608;
        15'h0802: data = 12'h607;
        15'h0803: data = 12'h600;
        15'h0804: data = 12'h602;
        15'h0805: data = 12'h603;
        15'h0806: data = 12'h604;
        15'h0807: data = 12'h605;
        15'h0808: data = 12'h60B;
        15'h0809: data = 12'h60C;
        15'h080A: data = 12'h60B;
        15'h080B: data = 12'h60B;
        15'h080C: data = 12'h600;
        15'h080D: data = 12'h605;
        15'h080E: data = 12'h600;
        15'h080F: data = 12'h5FF;
        15'h0810: data = 12'h607;
        15'h0811: data = 12'h608;
        15'h0812: data = 12'h60C;
        15'h0813: data = 12'h60E;
        15'h0814: data = 12'h60B;
        15'h0815: data = 12'h60C;
        15'h0816: data = 12'h605;
        15'h0817: data = 12'h601;
        15'h0818: data = 12'h5FD;
        15'h0819: data = 12'h604;
        15'h081A: data = 12'h607;
        15'h081B: data = 12'h62D;
        15'h081C: data = 12'h62C;
        15'h081D: data = 12'h629;
        15'h081E: data = 12'h62B;
        15'h081F: data = 12'h626;
        15'h0820: data = 12'h621;
        15'h0821: data = 12'h620;
        15'h0822: data = 12'h620;
        15'h0823: data = 12'h61E;
        15'h0824: data = 12'h625;
        15'h0825: data = 12'h629;
        15'h0826: data = 12'h62E;
        15'h0827: data = 12'h62A;
        15'h0828: data = 12'h628;
        15'h0829: data = 12'h625;
        15'h082A: data = 12'h61C;
        15'h082B: data = 12'h61E;
        15'h082C: data = 12'h61D;
        15'h082D: data = 12'h624;
        15'h082E: data = 12'h629;
        15'h082F: data = 12'h62B;
        15'h0830: data = 12'h62B;
        15'h0831: data = 12'h62A;
        15'h0832: data = 12'h626;
        15'h0833: data = 12'h620;
        15'h0834: data = 12'h61F;
        15'h0835: data = 12'h61F;
        15'h0836: data = 12'h624;
        15'h0837: data = 12'h627;
        15'h0838: data = 12'h628;
        15'h0839: data = 12'h62A;
        15'h083A: data = 12'h629;
        15'h083B: data = 12'h628;
        15'h083C: data = 12'h621;
        15'h083D: data = 12'h620;
        15'h083E: data = 12'h61F;
        15'h083F: data = 12'h61F;
        15'h0840: data = 12'h621;
        15'h0841: data = 12'h627;
        15'h0842: data = 12'h62A;
        15'h0843: data = 12'h62B;
        15'h0844: data = 12'h62A;
        15'h0845: data = 12'h626;
        15'h0846: data = 12'h625;
        15'h0847: data = 12'h620;
        15'h0848: data = 12'h61F;
        15'h0849: data = 12'h620;
        15'h084A: data = 12'h625;
        15'h084B: data = 12'h629;
        15'h084C: data = 12'h62B;
        15'h084D: data = 12'h62C;
        15'h084E: data = 12'h628;
        15'h084F: data = 12'h625;
        15'h0850: data = 12'h622;
        15'h0851: data = 12'h620;
        15'h0852: data = 12'h621;
        15'h0853: data = 12'h624;
        15'h0854: data = 12'h624;
        15'h0855: data = 12'h629;
        15'h0856: data = 12'h627;
        15'h0857: data = 12'h62C;
        15'h0858: data = 12'h62B;
        15'h0859: data = 12'h627;
        15'h085A: data = 12'h61E;
        15'h085B: data = 12'h620;
        15'h085C: data = 12'h628;
        15'h085D: data = 12'h642;
        15'h085E: data = 12'h64A;
        15'h085F: data = 12'h64A;
        15'h0860: data = 12'h64C;
        15'h0861: data = 12'h64B;
        15'h0862: data = 12'h647;
        15'h0863: data = 12'h642;
        15'h0864: data = 12'h640;
        15'h0865: data = 12'h63E;
        15'h0866: data = 12'h63F;
        15'h0867: data = 12'h641;
        15'h0868: data = 12'h647;
        15'h0869: data = 12'h64A;
        15'h086A: data = 12'h64A;
        15'h086B: data = 12'h649;
        15'h086C: data = 12'h646;
        15'h086D: data = 12'h63F;
        15'h086E: data = 12'h63E;
        15'h086F: data = 12'h63D;
        15'h0870: data = 12'h641;
        15'h0871: data = 12'h643;
        15'h0872: data = 12'h64A;
        15'h0873: data = 12'h64C;
        15'h0874: data = 12'h64D;
        15'h0875: data = 12'h647;
        15'h0876: data = 12'h643;
        15'h0877: data = 12'h63D;
        15'h0878: data = 12'h63B;
        15'h0879: data = 12'h63E;
        15'h087A: data = 12'h641;
        15'h087B: data = 12'h646;
        15'h087C: data = 12'h64C;
        15'h087D: data = 12'h64E;
        15'h087E: data = 12'h64B;
        15'h087F: data = 12'h647;
        15'h0880: data = 12'h641;
        15'h0881: data = 12'h63D;
        15'h0882: data = 12'h63F;
        15'h0883: data = 12'h63F;
        15'h0884: data = 12'h644;
        15'h0885: data = 12'h648;
        15'h0886: data = 12'h64C;
        15'h0887: data = 12'h64F;
        15'h0888: data = 12'h650;
        15'h0889: data = 12'h646;
        15'h088A: data = 12'h640;
        15'h088B: data = 12'h63A;
        15'h088C: data = 12'h63E;
        15'h088D: data = 12'h641;
        15'h088E: data = 12'h649;
        15'h088F: data = 12'h64A;
        15'h0890: data = 12'h64D;
        15'h0891: data = 12'h64B;
        15'h0892: data = 12'h649;
        15'h0893: data = 12'h647;
        15'h0894: data = 12'h641;
        15'h0895: data = 12'h640;
        15'h0896: data = 12'h640;
        15'h0897: data = 12'h643;
        15'h0898: data = 12'h647;
        15'h0899: data = 12'h64D;
        15'h089A: data = 12'h64D;
        15'h089B: data = 12'h64D;
        15'h089C: data = 12'h647;
        15'h089D: data = 12'h646;
        15'h089E: data = 12'h640;
        15'h089F: data = 12'h63C;
        15'h08A0: data = 12'h642;
        15'h08A1: data = 12'h644;
        15'h08A2: data = 12'h649;
        15'h08A3: data = 12'h64B;
        15'h08A4: data = 12'h64A;
        15'h08A5: data = 12'h647;
        15'h08A6: data = 12'h643;
        15'h08A7: data = 12'h642;
        15'h08A8: data = 12'h640;
        15'h08A9: data = 12'h63F;
        15'h08AA: data = 12'h646;
        15'h08AB: data = 12'h669;
        15'h08AC: data = 12'h66B;
        15'h08AD: data = 12'h66B;
        15'h08AE: data = 12'h66B;
        15'h08AF: data = 12'h66C;
        15'h08B0: data = 12'h667;
        15'h08B1: data = 12'h664;
        15'h08B2: data = 12'h662;
        15'h08B3: data = 12'h661;
        15'h08B4: data = 12'h661;
        15'h08B5: data = 12'h669;
        15'h08B6: data = 12'h66C;
        15'h08B7: data = 12'h66F;
        15'h08B8: data = 12'h66C;
        15'h08B9: data = 12'h666;
        15'h08BA: data = 12'h663;
        15'h08BB: data = 12'h664;
        15'h08BC: data = 12'h664;
        15'h08BD: data = 12'h665;
        15'h08BE: data = 12'h665;
        15'h08BF: data = 12'h66D;
        15'h08C0: data = 12'h66B;
        15'h08C1: data = 12'h66B;
        15'h08C2: data = 12'h66D;
        15'h08C3: data = 12'h667;
        15'h08C4: data = 12'h666;
        15'h08C5: data = 12'h665;
        15'h08C6: data = 12'h663;
        15'h08C7: data = 12'h664;
        15'h08C8: data = 12'h664;
        15'h08C9: data = 12'h66A;
        15'h08CA: data = 12'h66B;
        15'h08CB: data = 12'h66B;
        15'h08CC: data = 12'h66C;
        15'h08CD: data = 12'h66B;
        15'h08CE: data = 12'h662;
        15'h08CF: data = 12'h665;
        15'h08D0: data = 12'h663;
        15'h08D1: data = 12'h662;
        15'h08D2: data = 12'h667;
        15'h08D3: data = 12'h66C;
        15'h08D4: data = 12'h66F;
        15'h08D5: data = 12'h66B;
        15'h08D6: data = 12'h668;
        15'h08D7: data = 12'h666;
        15'h08D8: data = 12'h661;
        15'h08D9: data = 12'h65F;
        15'h08DA: data = 12'h65E;
        15'h08DB: data = 12'h662;
        15'h08DC: data = 12'h668;
        15'h08DD: data = 12'h66F;
        15'h08DE: data = 12'h670;
        15'h08DF: data = 12'h66C;
        15'h08E0: data = 12'h667;
        15'h08E1: data = 12'h660;
        15'h08E2: data = 12'h65E;
        15'h08E3: data = 12'h65E;
        15'h08E4: data = 12'h660;
        15'h08E5: data = 12'h664;
        15'h08E6: data = 12'h669;
        15'h08E7: data = 12'h66C;
        15'h08E8: data = 12'h66D;
        15'h08E9: data = 12'h66A;
        15'h08EA: data = 12'h665;
        15'h08EB: data = 12'h661;
        15'h08EC: data = 12'h65D;
        15'h08ED: data = 12'h661;
        15'h08EE: data = 12'h663;
        15'h08EF: data = 12'h667;
        15'h08F0: data = 12'h66E;
        15'h08F1: data = 12'h66B;
        15'h08F2: data = 12'h66D;
        15'h08F3: data = 12'h66A;
        15'h08F4: data = 12'h669;
        15'h08F5: data = 12'h663;
        15'h08F6: data = 12'h662;
        15'h08F7: data = 12'h665;
        15'h08F8: data = 12'h663;
        15'h08F9: data = 12'h668;
        15'h08FA: data = 12'h688;
        15'h08FB: data = 12'h68E;
        15'h08FC: data = 12'h68A;
        15'h08FD: data = 12'h685;
        15'h08FE: data = 12'h681;
        15'h08FF: data = 12'h683;
        15'h0900: data = 12'h67F;
        15'h0901: data = 12'h680;
        15'h0902: data = 12'h689;
        15'h0903: data = 12'h68A;
        15'h0904: data = 12'h68A;
        15'h0905: data = 12'h68B;
        15'h0906: data = 12'h68B;
        15'h0907: data = 12'h687;
        15'h0908: data = 12'h685;
        15'h0909: data = 12'h67E;
        15'h090A: data = 12'h67F;
        15'h090B: data = 12'h680;
        15'h090C: data = 12'h683;
        15'h090D: data = 12'h687;
        15'h090E: data = 12'h68B;
        15'h090F: data = 12'h68C;
        15'h0910: data = 12'h68B;
        15'h0911: data = 12'h686;
        15'h0912: data = 12'h680;
        15'h0913: data = 12'h67E;
        15'h0914: data = 12'h67E;
        15'h0915: data = 12'h682;
        15'h0916: data = 12'h687;
        15'h0917: data = 12'h68C;
        15'h0918: data = 12'h68C;
        15'h0919: data = 12'h689;
        15'h091A: data = 12'h687;
        15'h091B: data = 12'h682;
        15'h091C: data = 12'h67F;
        15'h091D: data = 12'h682;
        15'h091E: data = 12'h681;
        15'h091F: data = 12'h683;
        15'h0920: data = 12'h68A;
        15'h0921: data = 12'h68B;
        15'h0922: data = 12'h68A;
        15'h0923: data = 12'h688;
        15'h0924: data = 12'h683;
        15'h0925: data = 12'h681;
        15'h0926: data = 12'h680;
        15'h0927: data = 12'h67B;
        15'h0928: data = 12'h67F;
        15'h0929: data = 12'h687;
        15'h092A: data = 12'h686;
        15'h092B: data = 12'h689;
        15'h092C: data = 12'h68F;
        15'h092D: data = 12'h68B;
        15'h092E: data = 12'h687;
        15'h092F: data = 12'h683;
        15'h0930: data = 12'h682;
        15'h0931: data = 12'h67E;
        15'h0932: data = 12'h67E;
        15'h0933: data = 12'h682;
        15'h0934: data = 12'h688;
        15'h0935: data = 12'h68C;
        15'h0936: data = 12'h68F;
        15'h0937: data = 12'h689;
        15'h0938: data = 12'h681;
        15'h0939: data = 12'h682;
        15'h093A: data = 12'h67E;
        15'h093B: data = 12'h67F;
        15'h093C: data = 12'h683;
        15'h093D: data = 12'h687;
        15'h093E: data = 12'h68A;
        15'h093F: data = 12'h68E;
        15'h0940: data = 12'h68D;
        15'h0941: data = 12'h687;
        15'h0942: data = 12'h683;
        15'h0943: data = 12'h67E;
        15'h0944: data = 12'h681;
        15'h0945: data = 12'h67D;
        15'h0946: data = 12'h681;
        15'h0947: data = 12'h688;
        15'h0948: data = 12'h6A8;
        15'h0949: data = 12'h6A9;
        15'h094A: data = 12'h6A6;
        15'h094B: data = 12'h6A1;
        15'h094C: data = 12'h6A0;
        15'h094D: data = 12'h69C;
        15'h094E: data = 12'h69E;
        15'h094F: data = 12'h6A1;
        15'h0950: data = 12'h6A5;
        15'h0951: data = 12'h6AA;
        15'h0952: data = 12'h6A9;
        15'h0953: data = 12'h6A9;
        15'h0954: data = 12'h6A7;
        15'h0955: data = 12'h69E;
        15'h0956: data = 12'h6A1;
        15'h0957: data = 12'h69F;
        15'h0958: data = 12'h6A5;
        15'h0959: data = 12'h6A4;
        15'h095A: data = 12'h6A8;
        15'h095B: data = 12'h6A8;
        15'h095C: data = 12'h6A9;
        15'h095D: data = 12'h6AA;
        15'h095E: data = 12'h6A4;
        15'h095F: data = 12'h6A1;
        15'h0960: data = 12'h69F;
        15'h0961: data = 12'h6A0;
        15'h0962: data = 12'h6A1;
        15'h0963: data = 12'h6A2;
        15'h0964: data = 12'h6AC;
        15'h0965: data = 12'h6A8;
        15'h0966: data = 12'h6AB;
        15'h0967: data = 12'h6AD;
        15'h0968: data = 12'h6A9;
        15'h0969: data = 12'h6A3;
        15'h096A: data = 12'h69E;
        15'h096B: data = 12'h69C;
        15'h096C: data = 12'h6A1;
        15'h096D: data = 12'h6A6;
        15'h096E: data = 12'h6A7;
        15'h096F: data = 12'h6A7;
        15'h0970: data = 12'h6A9;
        15'h0971: data = 12'h6A7;
        15'h0972: data = 12'h6A4;
        15'h0973: data = 12'h6A2;
        15'h0974: data = 12'h6A0;
        15'h0975: data = 12'h6A0;
        15'h0976: data = 12'h6A1;
        15'h0977: data = 12'h6A6;
        15'h0978: data = 12'h6A7;
        15'h0979: data = 12'h6A9;
        15'h097A: data = 12'h6A8;
        15'h097B: data = 12'h6A5;
        15'h097C: data = 12'h6A5;
        15'h097D: data = 12'h6A3;
        15'h097E: data = 12'h6A2;
        15'h097F: data = 12'h69E;
        15'h0980: data = 12'h6A5;
        15'h0981: data = 12'h6A8;
        15'h0982: data = 12'h6A9;
        15'h0983: data = 12'h6AE;
        15'h0984: data = 12'h6AA;
        15'h0985: data = 12'h6A6;
        15'h0986: data = 12'h6A2;
        15'h0987: data = 12'h69F;
        15'h0988: data = 12'h69C;
        15'h0989: data = 12'h6A2;
        15'h098A: data = 12'h6A5;
        15'h098B: data = 12'h6AA;
        15'h098C: data = 12'h6AA;
        15'h098D: data = 12'h6AB;
        15'h098E: data = 12'h6AB;
        15'h098F: data = 12'h6A4;
        15'h0990: data = 12'h6A0;
        15'h0991: data = 12'h69D;
        15'h0992: data = 12'h69E;
        15'h0993: data = 12'h6A4;
        15'h0994: data = 12'h6AA;
        15'h0995: data = 12'h6B0;
        15'h0996: data = 12'h6A8;
        15'h0997: data = 12'h6C9;
        15'h0998: data = 12'h6C9;
        15'h0999: data = 12'h6C2;
        15'h099A: data = 12'h6BF;
        15'h099B: data = 12'h6BE;
        15'h099C: data = 12'h6C3;
        15'h099D: data = 12'h6C5;
        15'h099E: data = 12'h6C9;
        15'h099F: data = 12'h6CC;
        15'h09A0: data = 12'h6CA;
        15'h09A1: data = 12'h6CA;
        15'h09A2: data = 12'h6C5;
        15'h09A3: data = 12'h6C3;
        15'h09A4: data = 12'h6C3;
        15'h09A5: data = 12'h6BF;
        15'h09A6: data = 12'h6C5;
        15'h09A7: data = 12'h6CB;
        15'h09A8: data = 12'h6CB;
        15'h09A9: data = 12'h6CE;
        15'h09AA: data = 12'h6CE;
        15'h09AB: data = 12'h6CD;
        15'h09AC: data = 12'h6C4;
        15'h09AD: data = 12'h6C1;
        15'h09AE: data = 12'h6BF;
        15'h09AF: data = 12'h6C4;
        15'h09B0: data = 12'h6C6;
        15'h09B1: data = 12'h6C8;
        15'h09B2: data = 12'h6CF;
        15'h09B3: data = 12'h6CB;
        15'h09B4: data = 12'h6CB;
        15'h09B5: data = 12'h6C7;
        15'h09B6: data = 12'h6C1;
        15'h09B7: data = 12'h6BE;
        15'h09B8: data = 12'h6C0;
        15'h09B9: data = 12'h6C3;
        15'h09BA: data = 12'h6C5;
        15'h09BB: data = 12'h6CD;
        15'h09BC: data = 12'h6C9;
        15'h09BD: data = 12'h6C9;
        15'h09BE: data = 12'h6C9;
        15'h09BF: data = 12'h6BE;
        15'h09C0: data = 12'h6BB;
        15'h09C1: data = 12'h6BE;
        15'h09C2: data = 12'h6BE;
        15'h09C3: data = 12'h6C3;
        15'h09C4: data = 12'h6C7;
        15'h09C5: data = 12'h6CB;
        15'h09C6: data = 12'h6C7;
        15'h09C7: data = 12'h6C8;
        15'h09C8: data = 12'h6C7;
        15'h09C9: data = 12'h6BF;
        15'h09CA: data = 12'h6C0;
        15'h09CB: data = 12'h6BE;
        15'h09CC: data = 12'h6C0;
        15'h09CD: data = 12'h6C6;
        15'h09CE: data = 12'h6C7;
        15'h09CF: data = 12'h6CB;
        15'h09D0: data = 12'h6C9;
        15'h09D1: data = 12'h6C6;
        15'h09D2: data = 12'h6C3;
        15'h09D3: data = 12'h6C1;
        15'h09D4: data = 12'h6BD;
        15'h09D5: data = 12'h6BD;
        15'h09D6: data = 12'h6C0;
        15'h09D7: data = 12'h6C8;
        15'h09D8: data = 12'h6C7;
        15'h09D9: data = 12'h6CC;
        15'h09DA: data = 12'h6CC;
        15'h09DB: data = 12'h6C9;
        15'h09DC: data = 12'h6C5;
        15'h09DD: data = 12'h6BE;
        15'h09DE: data = 12'h6C1;
        15'h09DF: data = 12'h6C4;
        15'h09E0: data = 12'h6C7;
        15'h09E1: data = 12'h6C8;
        15'h09E2: data = 12'h6C9;
        15'h09E3: data = 12'h6CB;
        15'h09E4: data = 12'h6C6;
        15'h09E5: data = 12'h6C1;
        15'h09E6: data = 12'h6BE;
        15'h09E7: data = 12'h6BE;
        15'h09E8: data = 12'h6BE;
        15'h09E9: data = 12'h6C1;
        15'h09EA: data = 12'h6CA;
        15'h09EB: data = 12'h6C8;
        15'h09EC: data = 12'h6CB;
        15'h09ED: data = 12'h6C9;
        15'h09EE: data = 12'h6C9;
        15'h09EF: data = 12'h6C5;
        15'h09F0: data = 12'h6BF;
        15'h09F1: data = 12'h6BE;
        15'h09F2: data = 12'h6C0;
        15'h09F3: data = 12'h6DE;
        15'h09F4: data = 12'h6E7;
        15'h09F5: data = 12'h6E7;
        15'h09F6: data = 12'h6EA;
        15'h09F7: data = 12'h6EC;
        15'h09F8: data = 12'h6E7;
        15'h09F9: data = 12'h6E1;
        15'h09FA: data = 12'h6DF;
        15'h09FB: data = 12'h6DD;
        15'h09FC: data = 12'h6E0;
        15'h09FD: data = 12'h6E6;
        15'h09FE: data = 12'h6E8;
        15'h09FF: data = 12'h6EE;
        15'h0A00: data = 12'h6EF;
        15'h0A01: data = 12'h6EB;
        15'h0A02: data = 12'h6E5;
        15'h0A03: data = 12'h6E0;
        15'h0A04: data = 12'h6E0;
        15'h0A05: data = 12'h6DE;
        15'h0A06: data = 12'h6E1;
        15'h0A07: data = 12'h6E8;
        15'h0A08: data = 12'h6EC;
        15'h0A09: data = 12'h6F0;
        15'h0A0A: data = 12'h6EC;
        15'h0A0B: data = 12'h6EB;
        15'h0A0C: data = 12'h6E5;
        15'h0A0D: data = 12'h6E0;
        15'h0A0E: data = 12'h6DC;
        15'h0A0F: data = 12'h6DC;
        15'h0A10: data = 12'h6E2;
        15'h0A11: data = 12'h6EB;
        15'h0A12: data = 12'h6EE;
        15'h0A13: data = 12'h6EA;
        15'h0A14: data = 12'h6EB;
        15'h0A15: data = 12'h6E3;
        15'h0A16: data = 12'h6DE;
        15'h0A17: data = 12'h6E1;
        15'h0A18: data = 12'h6DC;
        15'h0A19: data = 12'h6E0;
        15'h0A1A: data = 12'h6E3;
        15'h0A1B: data = 12'h6E9;
        15'h0A1C: data = 12'h6ED;
        15'h0A1D: data = 12'h6E8;
        15'h0A1E: data = 12'h6E8;
        15'h0A1F: data = 12'h6DF;
        15'h0A20: data = 12'h6DF;
        15'h0A21: data = 12'h6DD;
        15'h0A22: data = 12'h6DE;
        15'h0A23: data = 12'h6E1;
        15'h0A24: data = 12'h6E8;
        15'h0A25: data = 12'h6E9;
        15'h0A26: data = 12'h6E9;
        15'h0A27: data = 12'h6EA;
        15'h0A28: data = 12'h6E5;
        15'h0A29: data = 12'h6E4;
        15'h0A2A: data = 12'h6E1;
        15'h0A2B: data = 12'h6DE;
        15'h0A2C: data = 12'h6DF;
        15'h0A2D: data = 12'h6E4;
        15'h0A2E: data = 12'h6E7;
        15'h0A2F: data = 12'h6EA;
        15'h0A30: data = 12'h6EA;
        15'h0A31: data = 12'h6EC;
        15'h0A32: data = 12'h6E5;
        15'h0A33: data = 12'h6E2;
        15'h0A34: data = 12'h6FE;
        15'h0A35: data = 12'h6FC;
        15'h0A36: data = 12'h702;
        15'h0A37: data = 12'h708;
        15'h0A38: data = 12'h707;
        15'h0A39: data = 12'h70C;
        15'h0A3A: data = 12'h70A;
        15'h0A3B: data = 12'h709;
        15'h0A3C: data = 12'h700;
        15'h0A3D: data = 12'h6FC;
        15'h0A3E: data = 12'h6FC;
        15'h0A3F: data = 12'h701;
        15'h0A40: data = 12'h704;
        15'h0A41: data = 12'h706;
        15'h0A42: data = 12'h705;
        15'h0A43: data = 12'h707;
        15'h0A44: data = 12'h70B;
        15'h0A45: data = 12'h707;
        15'h0A46: data = 12'h701;
        15'h0A47: data = 12'h6FE;
        15'h0A48: data = 12'h6FF;
        15'h0A49: data = 12'h6FF;
        15'h0A4A: data = 12'h704;
        15'h0A4B: data = 12'h705;
        15'h0A4C: data = 12'h70B;
        15'h0A4D: data = 12'h709;
        15'h0A4E: data = 12'h707;
        15'h0A4F: data = 12'h703;
        15'h0A50: data = 12'h6FE;
        15'h0A51: data = 12'h6FF;
        15'h0A52: data = 12'h6FD;
        15'h0A53: data = 12'h6FE;
        15'h0A54: data = 12'h702;
        15'h0A55: data = 12'h709;
        15'h0A56: data = 12'h709;
        15'h0A57: data = 12'h707;
        15'h0A58: data = 12'h705;
        15'h0A59: data = 12'h6FF;
        15'h0A5A: data = 12'h6FD;
        15'h0A5B: data = 12'h6FF;
        15'h0A5C: data = 12'h6FC;
        15'h0A5D: data = 12'h702;
        15'h0A5E: data = 12'h707;
        15'h0A5F: data = 12'h70B;
        15'h0A60: data = 12'h706;
        15'h0A61: data = 12'h708;
        15'h0A62: data = 12'h700;
        15'h0A63: data = 12'h6FE;
        15'h0A64: data = 12'h6FE;
        15'h0A65: data = 12'h701;
        15'h0A66: data = 12'h700;
        15'h0A67: data = 12'h70A;
        15'h0A68: data = 12'h706;
        15'h0A69: data = 12'h70B;
        15'h0A6A: data = 12'h709;
        15'h0A6B: data = 12'h706;
        15'h0A6C: data = 12'h700;
        15'h0A6D: data = 12'h6FD;
        15'h0A6E: data = 12'h6FB;
        15'h0A6F: data = 12'h6FB;
        15'h0A70: data = 12'h701;
        15'h0A71: data = 12'h705;
        15'h0A72: data = 12'h705;
        15'h0A73: data = 12'h707;
        15'h0A74: data = 12'h707;
        15'h0A75: data = 12'h707;
        15'h0A76: data = 12'h704;
        15'h0A77: data = 12'h700;
        15'h0A78: data = 12'h6FF;
        15'h0A79: data = 12'h6FD;
        15'h0A7A: data = 12'h701;
        15'h0A7B: data = 12'h703;
        15'h0A7C: data = 12'h70B;
        15'h0A7D: data = 12'h70C;
        15'h0A7E: data = 12'h70A;
        15'h0A7F: data = 12'h706;
        15'h0A80: data = 12'h702;
        15'h0A81: data = 12'h6FE;
        15'h0A82: data = 12'h6FF;
        15'h0A83: data = 12'h719;
        15'h0A84: data = 12'h718;
        15'h0A85: data = 12'h71E;
        15'h0A86: data = 12'h720;
        15'h0A87: data = 12'h720;
        15'h0A88: data = 12'h71F;
        15'h0A89: data = 12'h718;
        15'h0A8A: data = 12'h714;
        15'h0A8B: data = 12'h716;
        15'h0A8C: data = 12'h716;
        15'h0A8D: data = 12'h71C;
        15'h0A8E: data = 12'h71C;
        15'h0A8F: data = 12'h724;
        15'h0A90: data = 12'h724;
        15'h0A91: data = 12'h71F;
        15'h0A92: data = 12'h71F;
        15'h0A93: data = 12'h716;
        15'h0A94: data = 12'h712;
        15'h0A95: data = 12'h713;
        15'h0A96: data = 12'h716;
        15'h0A97: data = 12'h71A;
        15'h0A98: data = 12'h723;
        15'h0A99: data = 12'h724;
        15'h0A9A: data = 12'h71F;
        15'h0A9B: data = 12'h71E;
        15'h0A9C: data = 12'h71A;
        15'h0A9D: data = 12'h715;
        15'h0A9E: data = 12'h714;
        15'h0A9F: data = 12'h716;
        15'h0AA0: data = 12'h71A;
        15'h0AA1: data = 12'h71E;
        15'h0AA2: data = 12'h71F;
        15'h0AA3: data = 12'h722;
        15'h0AA4: data = 12'h71F;
        15'h0AA5: data = 12'h71B;
        15'h0AA6: data = 12'h719;
        15'h0AA7: data = 12'h711;
        15'h0AA8: data = 12'h715;
        15'h0AA9: data = 12'h716;
        15'h0AAA: data = 12'h71C;
        15'h0AAB: data = 12'h720;
        15'h0AAC: data = 12'h722;
        15'h0AAD: data = 12'h722;
        15'h0AAE: data = 12'h71E;
        15'h0AAF: data = 12'h71D;
        15'h0AB0: data = 12'h719;
        15'h0AB1: data = 12'h718;
        15'h0AB2: data = 12'h716;
        15'h0AB3: data = 12'h71A;
        15'h0AB4: data = 12'h71E;
        15'h0AB5: data = 12'h71F;
        15'h0AB6: data = 12'h71D;
        15'h0AB7: data = 12'h71E;
        15'h0AB8: data = 12'h71D;
        15'h0AB9: data = 12'h719;
        15'h0ABA: data = 12'h715;
        15'h0ABB: data = 12'h714;
        15'h0ABC: data = 12'h713;
        15'h0ABD: data = 12'h717;
        15'h0ABE: data = 12'h71E;
        15'h0ABF: data = 12'h721;
        15'h0AC0: data = 12'h71F;
        15'h0AC1: data = 12'h723;
        15'h0AC2: data = 12'h71A;
        15'h0AC3: data = 12'h719;
        15'h0AC4: data = 12'h713;
        15'h0AC5: data = 12'h716;
        15'h0AC6: data = 12'h718;
        15'h0AC7: data = 12'h71D;
        15'h0AC8: data = 12'h71E;
        15'h0AC9: data = 12'h721;
        15'h0ACA: data = 12'h722;
        15'h0ACB: data = 12'h722;
        15'h0ACC: data = 12'h71C;
        15'h0ACD: data = 12'h718;
        15'h0ACE: data = 12'h713;
        15'h0ACF: data = 12'h714;
        15'h0AD0: data = 12'h718;
        15'h0AD1: data = 12'h71E;
        15'h0AD2: data = 12'h73F;
        15'h0AD3: data = 12'h741;
        15'h0AD4: data = 12'h73F;
        15'h0AD5: data = 12'h73C;
        15'h0AD6: data = 12'h736;
        15'h0AD7: data = 12'h736;
        15'h0AD8: data = 12'h732;
        15'h0AD9: data = 12'h735;
        15'h0ADA: data = 12'h73B;
        15'h0ADB: data = 12'h73F;
        15'h0ADC: data = 12'h741;
        15'h0ADD: data = 12'h744;
        15'h0ADE: data = 12'h73F;
        15'h0ADF: data = 12'h73A;
        15'h0AE0: data = 12'h735;
        15'h0AE1: data = 12'h734;
        15'h0AE2: data = 12'h736;
        15'h0AE3: data = 12'h739;
        15'h0AE4: data = 12'h73F;
        15'h0AE5: data = 12'h741;
        15'h0AE6: data = 12'h745;
        15'h0AE7: data = 12'h743;
        15'h0AE8: data = 12'h73F;
        15'h0AE9: data = 12'h73D;
        15'h0AEA: data = 12'h73B;
        15'h0AEB: data = 12'h735;
        15'h0AEC: data = 12'h736;
        15'h0AED: data = 12'h73B;
        15'h0AEE: data = 12'h73D;
        15'h0AEF: data = 12'h73E;
        15'h0AF0: data = 12'h73D;
        15'h0AF1: data = 12'h742;
        15'h0AF2: data = 12'h73E;
        15'h0AF3: data = 12'h737;
        15'h0AF4: data = 12'h737;
        15'h0AF5: data = 12'h736;
        15'h0AF6: data = 12'h736;
        15'h0AF7: data = 12'h73F;
        15'h0AF8: data = 12'h741;
        15'h0AF9: data = 12'h741;
        15'h0AFA: data = 12'h740;
        15'h0AFB: data = 12'h73F;
        15'h0AFC: data = 12'h73C;
        15'h0AFD: data = 12'h738;
        15'h0AFE: data = 12'h736;
        15'h0AFF: data = 12'h735;
        15'h0B00: data = 12'h734;
        15'h0B01: data = 12'h73B;
        15'h0B02: data = 12'h73E;
        15'h0B03: data = 12'h741;
        15'h0B04: data = 12'h744;
        15'h0B05: data = 12'h741;
        15'h0B06: data = 12'h73B;
        15'h0B07: data = 12'h735;
        15'h0B08: data = 12'h732;
        15'h0B09: data = 12'h734;
        15'h0B0A: data = 12'h738;
        15'h0B0B: data = 12'h740;
        15'h0B0C: data = 12'h741;
        15'h0B0D: data = 12'h744;
        15'h0B0E: data = 12'h740;
        15'h0B0F: data = 12'h743;
        15'h0B10: data = 12'h73C;
        15'h0B11: data = 12'h738;
        15'h0B12: data = 12'h734;
        15'h0B13: data = 12'h75A;
        15'h0B14: data = 12'h75D;
        15'h0B15: data = 12'h760;
        15'h0B16: data = 12'h761;
        15'h0B17: data = 12'h761;
        15'h0B18: data = 12'h75F;
        15'h0B19: data = 12'h75A;
        15'h0B1A: data = 12'h755;
        15'h0B1B: data = 12'h755;
        15'h0B1C: data = 12'h754;
        15'h0B1D: data = 12'h758;
        15'h0B1E: data = 12'h75C;
        15'h0B1F: data = 12'h75F;
        15'h0B20: data = 12'h763;
        15'h0B21: data = 12'h763;
        15'h0B22: data = 12'h762;
        15'h0B23: data = 12'h759;
        15'h0B24: data = 12'h758;
        15'h0B25: data = 12'h757;
        15'h0B26: data = 12'h754;
        15'h0B27: data = 12'h757;
        15'h0B28: data = 12'h75D;
        15'h0B29: data = 12'h75E;
        15'h0B2A: data = 12'h762;
        15'h0B2B: data = 12'h75F;
        15'h0B2C: data = 12'h75B;
        15'h0B2D: data = 12'h758;
        15'h0B2E: data = 12'h759;
        15'h0B2F: data = 12'h758;
        15'h0B30: data = 12'h759;
        15'h0B31: data = 12'h75D;
        15'h0B32: data = 12'h763;
        15'h0B33: data = 12'h760;
        15'h0B34: data = 12'h761;
        15'h0B35: data = 12'h75F;
        15'h0B36: data = 12'h75B;
        15'h0B37: data = 12'h759;
        15'h0B38: data = 12'h757;
        15'h0B39: data = 12'h757;
        15'h0B3A: data = 12'h756;
        15'h0B3B: data = 12'h75A;
        15'h0B3C: data = 12'h75F;
        15'h0B3D: data = 12'h760;
        15'h0B3E: data = 12'h760;
        15'h0B3F: data = 12'h75F;
        15'h0B40: data = 12'h75C;
        15'h0B41: data = 12'h75A;
        15'h0B42: data = 12'h754;
        15'h0B43: data = 12'h753;
        15'h0B44: data = 12'h753;
        15'h0B45: data = 12'h75D;
        15'h0B46: data = 12'h761;
        15'h0B47: data = 12'h763;
        15'h0B48: data = 12'h760;
        15'h0B49: data = 12'h761;
        15'h0B4A: data = 12'h75B;
        15'h0B4B: data = 12'h756;
        15'h0B4C: data = 12'h755;
        15'h0B4D: data = 12'h753;
        15'h0B4E: data = 12'h758;
        15'h0B4F: data = 12'h75E;
        15'h0B50: data = 12'h763;
        15'h0B51: data = 12'h764;
        15'h0B52: data = 12'h766;
        15'h0B53: data = 12'h75C;
        15'h0B54: data = 12'h75A;
        15'h0B55: data = 12'h757;
        15'h0B56: data = 12'h754;
        15'h0B57: data = 12'h755;
        15'h0B58: data = 12'h75B;
        15'h0B59: data = 12'h761;
        15'h0B5A: data = 12'h762;
        15'h0B5B: data = 12'h764;
        15'h0B5C: data = 12'h761;
        15'h0B5D: data = 12'h75F;
        15'h0B5E: data = 12'h756;
        15'h0B5F: data = 12'h757;
        15'h0B60: data = 12'h758;
        15'h0B61: data = 12'h758;
        15'h0B62: data = 12'h75D;
        15'h0B63: data = 12'h760;
        15'h0B64: data = 12'h763;
        15'h0B65: data = 12'h75F;
        15'h0B66: data = 12'h762;
        15'h0B67: data = 12'h75D;
        15'h0B68: data = 12'h759;
        15'h0B69: data = 12'h758;
        15'h0B6A: data = 12'h757;
        15'h0B6B: data = 12'h756;
        15'h0B6C: data = 12'h75C;
        15'h0B6D: data = 12'h75B;
        15'h0B6E: data = 12'h75D;
        15'h0B6F: data = 12'h77E;
        15'h0B70: data = 12'h780;
        15'h0B71: data = 12'h77F;
        15'h0B72: data = 12'h77C;
        15'h0B73: data = 12'h777;
        15'h0B74: data = 12'h778;
        15'h0B75: data = 12'h778;
        15'h0B76: data = 12'h77D;
        15'h0B77: data = 12'h77D;
        15'h0B78: data = 12'h780;
        15'h0B79: data = 12'h782;
        15'h0B7A: data = 12'h782;
        15'h0B7B: data = 12'h77D;
        15'h0B7C: data = 12'h775;
        15'h0B7D: data = 12'h778;
        15'h0B7E: data = 12'h779;
        15'h0B7F: data = 12'h779;
        15'h0B80: data = 12'h77D;
        15'h0B81: data = 12'h785;
        15'h0B82: data = 12'h785;
        15'h0B83: data = 12'h783;
        15'h0B84: data = 12'h782;
        15'h0B85: data = 12'h77C;
        15'h0B86: data = 12'h777;
        15'h0B87: data = 12'h778;
        15'h0B88: data = 12'h776;
        15'h0B89: data = 12'h779;
        15'h0B8A: data = 12'h77C;
        15'h0B8B: data = 12'h784;
        15'h0B8C: data = 12'h781;
        15'h0B8D: data = 12'h783;
        15'h0B8E: data = 12'h77C;
        15'h0B8F: data = 12'h77A;
        15'h0B90: data = 12'h776;
        15'h0B91: data = 12'h778;
        15'h0B92: data = 12'h776;
        15'h0B93: data = 12'h778;
        15'h0B94: data = 12'h784;
        15'h0B95: data = 12'h782;
        15'h0B96: data = 12'h781;
        15'h0B97: data = 12'h784;
        15'h0B98: data = 12'h77B;
        15'h0B99: data = 12'h779;
        15'h0B9A: data = 12'h774;
        15'h0B9B: data = 12'h779;
        15'h0B9C: data = 12'h77A;
        15'h0B9D: data = 12'h781;
        15'h0B9E: data = 12'h784;
        15'h0B9F: data = 12'h784;
        15'h0BA0: data = 12'h77F;
        15'h0BA1: data = 12'h780;
        15'h0BA2: data = 12'h77D;
        15'h0BA3: data = 12'h77A;
        15'h0BA4: data = 12'h77A;
        15'h0BA5: data = 12'h776;
        15'h0BA6: data = 12'h77A;
        15'h0BA7: data = 12'h77C;
        15'h0BA8: data = 12'h77C;
        15'h0BA9: data = 12'h781;
        15'h0BAA: data = 12'h77F;
        15'h0BAB: data = 12'h77E;
        15'h0BAC: data = 12'h77C;
        15'h0BAD: data = 12'h778;
        15'h0BAE: data = 12'h777;
        15'h0BAF: data = 12'h779;
        15'h0BB0: data = 12'h792;
        15'h0BB1: data = 12'h79C;
        15'h0BB2: data = 12'h7A0;
        15'h0BB3: data = 12'h7A1;
        15'h0BB4: data = 12'h79E;
        15'h0BB5: data = 12'h79A;
        15'h0BB6: data = 12'h79A;
        15'h0BB7: data = 12'h796;
        15'h0BB8: data = 12'h79F;
        15'h0BB9: data = 12'h79C;
        15'h0BBA: data = 12'h79F;
        15'h0BBB: data = 12'h79D;
        15'h0BBC: data = 12'h7A2;
        15'h0BBD: data = 12'h7A0;
        15'h0BBE: data = 12'h79B;
        15'h0BBF: data = 12'h79E;
        15'h0BC0: data = 12'h79C;
        15'h0BC1: data = 12'h79D;
        15'h0BC2: data = 12'h798;
        15'h0BC3: data = 12'h79D;
        15'h0BC4: data = 12'h79D;
        15'h0BC5: data = 12'h7A3;
        15'h0BC6: data = 12'h7A3;
        15'h0BC7: data = 12'h7A2;
        15'h0BC8: data = 12'h79F;
        15'h0BC9: data = 12'h799;
        15'h0BCA: data = 12'h797;
        15'h0BCB: data = 12'h793;
        15'h0BCC: data = 12'h798;
        15'h0BCD: data = 12'h798;
        15'h0BCE: data = 12'h79C;
        15'h0BCF: data = 12'h79E;
        15'h0BD0: data = 12'h7A3;
        15'h0BD1: data = 12'h7A1;
        15'h0BD2: data = 12'h79D;
        15'h0BD3: data = 12'h79A;
        15'h0BD4: data = 12'h796;
        15'h0BD5: data = 12'h793;
        15'h0BD6: data = 12'h794;
        15'h0BD7: data = 12'h798;
        15'h0BD8: data = 12'h79F;
        15'h0BD9: data = 12'h7A3;
        15'h0BDA: data = 12'h79F;
        15'h0BDB: data = 12'h7A1;
        15'h0BDC: data = 12'h79E;
        15'h0BDD: data = 12'h799;
        15'h0BDE: data = 12'h797;
        15'h0BDF: data = 12'h793;
        15'h0BE0: data = 12'h797;
        15'h0BE1: data = 12'h79B;
        15'h0BE2: data = 12'h7A0;
        15'h0BE3: data = 12'h7A2;
        15'h0BE4: data = 12'h7A1;
        15'h0BE5: data = 12'h79E;
        15'h0BE6: data = 12'h79F;
        15'h0BE7: data = 12'h797;
        15'h0BE8: data = 12'h794;
        15'h0BE9: data = 12'h790;
        15'h0BEA: data = 12'h791;
        15'h0BEB: data = 12'h799;
        15'h0BEC: data = 12'h7A1;
        15'h0BED: data = 12'h7A3;
        15'h0BEE: data = 12'h7A0;
        15'h0BEF: data = 12'h7A1;
        15'h0BF0: data = 12'h79E;
        15'h0BF1: data = 12'h799;
        15'h0BF2: data = 12'h797;
        15'h0BF3: data = 12'h792;
        15'h0BF4: data = 12'h794;
        15'h0BF5: data = 12'h79B;
        15'h0BF6: data = 12'h79E;
        15'h0BF7: data = 12'h7A0;
        15'h0BF8: data = 12'h79F;
        15'h0BF9: data = 12'h79B;
        15'h0BFA: data = 12'h79A;
        15'h0BFB: data = 12'h79A;
        15'h0BFC: data = 12'h795;
        15'h0BFD: data = 12'h795;
        15'h0BFE: data = 12'h794;
        15'h0BFF: data = 12'h7BB;
        15'h0C00: data = 12'h7BC;
        15'h0C01: data = 12'h7C5;
        15'h0C02: data = 12'h7C1;
        15'h0C03: data = 12'h7C0;
        15'h0C04: data = 12'h7BA;
        15'h0C05: data = 12'h7B7;
        15'h0C06: data = 12'h7B5;
        15'h0C07: data = 12'h7B5;
        15'h0C08: data = 12'h7B8;
        15'h0C09: data = 12'h7BE;
        15'h0C0A: data = 12'h7BF;
        15'h0C0B: data = 12'h7C2;
        15'h0C0C: data = 12'h7BF;
        15'h0C0D: data = 12'h7BD;
        15'h0C0E: data = 12'h7C0;
        15'h0C0F: data = 12'h7B9;
        15'h0C10: data = 12'h7BA;
        15'h0C11: data = 12'h7B9;
        15'h0C12: data = 12'h7B8;
        15'h0C13: data = 12'h7BD;
        15'h0C14: data = 12'h7BF;
        15'h0C15: data = 12'h7C4;
        15'h0C16: data = 12'h7C0;
        15'h0C17: data = 12'h7C1;
        15'h0C18: data = 12'h7BE;
        15'h0C19: data = 12'h7BA;
        15'h0C1A: data = 12'h7B7;
        15'h0C1B: data = 12'h7B6;
        15'h0C1C: data = 12'h7B2;
        15'h0C1D: data = 12'h7BB;
        15'h0C1E: data = 12'h7C2;
        15'h0C1F: data = 12'h7C3;
        15'h0C20: data = 12'h7C4;
        15'h0C21: data = 12'h7C4;
        15'h0C22: data = 12'h7BB;
        15'h0C23: data = 12'h7BA;
        15'h0C24: data = 12'h7B3;
        15'h0C25: data = 12'h7B6;
        15'h0C26: data = 12'h7B7;
        15'h0C27: data = 12'h7BC;
        15'h0C28: data = 12'h7BE;
        15'h0C29: data = 12'h7C2;
        15'h0C2A: data = 12'h7C2;
        15'h0C2B: data = 12'h7BE;
        15'h0C2C: data = 12'h7BA;
        15'h0C2D: data = 12'h7B4;
        15'h0C2E: data = 12'h7B3;
        15'h0C2F: data = 12'h7B6;
        15'h0C30: data = 12'h7BB;
        15'h0C31: data = 12'h7BD;
        15'h0C32: data = 12'h7C0;
        15'h0C33: data = 12'h7C2;
        15'h0C34: data = 12'h7C0;
        15'h0C35: data = 12'h7C0;
        15'h0C36: data = 12'h7B7;
        15'h0C37: data = 12'h7B2;
        15'h0C38: data = 12'h7B9;
        15'h0C39: data = 12'h7B9;
        15'h0C3A: data = 12'h7BE;
        15'h0C3B: data = 12'h7C2;
        15'h0C3C: data = 12'h7C1;
        15'h0C3D: data = 12'h7C0;
        15'h0C3E: data = 12'h7BE;
        15'h0C3F: data = 12'h7BC;
        15'h0C40: data = 12'h7B6;
        15'h0C41: data = 12'h7CF;
        15'h0C42: data = 12'h7DB;
        15'h0C43: data = 12'h7DB;
        15'h0C44: data = 12'h7DD;
        15'h0C45: data = 12'h7E0;
        15'h0C46: data = 12'h7E2;
        15'h0C47: data = 12'h7DF;
        15'h0C48: data = 12'h7DD;
        15'h0C49: data = 12'h7DB;
        15'h0C4A: data = 12'h7D9;
        15'h0C4B: data = 12'h7D5;
        15'h0C4C: data = 12'h7D5;
        15'h0C4D: data = 12'h7DA;
        15'h0C4E: data = 12'h7DC;
        15'h0C4F: data = 12'h7E0;
        15'h0C50: data = 12'h7E3;
        15'h0C51: data = 12'h7E2;
        15'h0C52: data = 12'h7DE;
        15'h0C53: data = 12'h7DD;
        15'h0C54: data = 12'h7D6;
        15'h0C55: data = 12'h7CF;
        15'h0C56: data = 12'h7D4;
        15'h0C57: data = 12'h7D7;
        15'h0C58: data = 12'h7D9;
        15'h0C59: data = 12'h7DF;
        15'h0C5A: data = 12'h7E2;
        15'h0C5B: data = 12'h7DE;
        15'h0C5C: data = 12'h7DD;
        15'h0C5D: data = 12'h7DA;
        15'h0C5E: data = 12'h7D5;
        15'h0C5F: data = 12'h7D2;
        15'h0C60: data = 12'h7D3;
        15'h0C61: data = 12'h7D8;
        15'h0C62: data = 12'h7DD;
        15'h0C63: data = 12'h7E4;
        15'h0C64: data = 12'h7E2;
        15'h0C65: data = 12'h7E1;
        15'h0C66: data = 12'h7DF;
        15'h0C67: data = 12'h7D6;
        15'h0C68: data = 12'h7D1;
        15'h0C69: data = 12'h7D1;
        15'h0C6A: data = 12'h7D4;
        15'h0C6B: data = 12'h7D8;
        15'h0C6C: data = 12'h7DF;
        15'h0C6D: data = 12'h7DF;
        15'h0C6E: data = 12'h7E1;
        15'h0C6F: data = 12'h7E1;
        15'h0C70: data = 12'h7E2;
        15'h0C71: data = 12'h7D9;
        15'h0C72: data = 12'h7DA;
        15'h0C73: data = 12'h7D6;
        15'h0C74: data = 12'h7D3;
        15'h0C75: data = 12'h7DB;
        15'h0C76: data = 12'h7DF;
        15'h0C77: data = 12'h7E1;
        15'h0C78: data = 12'h7E1;
        15'h0C79: data = 12'h7E4;
        15'h0C7A: data = 12'h7DF;
        15'h0C7B: data = 12'h7D7;
        15'h0C7C: data = 12'h7D2;
        15'h0C7D: data = 12'h7D3;
        15'h0C7E: data = 12'h7D6;
        15'h0C7F: data = 12'h7DF;
        15'h0C80: data = 12'h7E1;
        15'h0C81: data = 12'h7E4;
        15'h0C82: data = 12'h7E3;
        15'h0C83: data = 12'h7E1;
        15'h0C84: data = 12'h7DF;
        15'h0C85: data = 12'h7D9;
        15'h0C86: data = 12'h7D6;
        15'h0C87: data = 12'h7D5;
        15'h0C88: data = 12'h7D8;
        15'h0C89: data = 12'h7DD;
        15'h0C8A: data = 12'h7E0;
        15'h0C8B: data = 12'h7E0;
        15'h0C8C: data = 12'h7E3;
        15'h0C8D: data = 12'h7E1;
        15'h0C8E: data = 12'h7DF;
        15'h0C8F: data = 12'h7F9;
        15'h0C90: data = 12'h7F2;
        15'h0C91: data = 12'h7F4;
        15'h0C92: data = 12'h7FA;
        15'h0C93: data = 12'h7FC;
        15'h0C94: data = 12'h7FB;
        15'h0C95: data = 12'h804;
        15'h0C96: data = 12'h803;
        15'h0C97: data = 12'h803;
        15'h0C98: data = 12'h7FD;
        15'h0C99: data = 12'h7F7;
        15'h0C9A: data = 12'h7F8;
        15'h0C9B: data = 12'h7F8;
        15'h0C9C: data = 12'h7F5;
        15'h0C9D: data = 12'h7FB;
        15'h0C9E: data = 12'h800;
        15'h0C9F: data = 12'h802;
        15'h0CA0: data = 12'h802;
        15'h0CA1: data = 12'h802;
        15'h0CA2: data = 12'h7FD;
        15'h0CA3: data = 12'h7F8;
        15'h0CA4: data = 12'h7F6;
        15'h0CA5: data = 12'h7F3;
        15'h0CA6: data = 12'h7F9;
        15'h0CA7: data = 12'h7FB;
        15'h0CA8: data = 12'h800;
        15'h0CA9: data = 12'h804;
        15'h0CAA: data = 12'h805;
        15'h0CAB: data = 12'h804;
        15'h0CAC: data = 12'h7FD;
        15'h0CAD: data = 12'h7F7;
        15'h0CAE: data = 12'h7F6;
        15'h0CAF: data = 12'h7F3;
        15'h0CB0: data = 12'h7F6;
        15'h0CB1: data = 12'h7FD;
        15'h0CB2: data = 12'h805;
        15'h0CB3: data = 12'h802;
        15'h0CB4: data = 12'h804;
        15'h0CB5: data = 12'h7FF;
        15'h0CB6: data = 12'h7FA;
        15'h0CB7: data = 12'h7F5;
        15'h0CB8: data = 12'h7F5;
        15'h0CB9: data = 12'h7F6;
        15'h0CBA: data = 12'h7FB;
        15'h0CBB: data = 12'h7FC;
        15'h0CBC: data = 12'h7FD;
        15'h0CBD: data = 12'h7FF;
        15'h0CBE: data = 12'h7FF;
        15'h0CBF: data = 12'h7FF;
        15'h0CC0: data = 12'h7FB;
        15'h0CC1: data = 12'h7F8;
        15'h0CC2: data = 12'h7F6;
        15'h0CC3: data = 12'h7F5;
        15'h0CC4: data = 12'h7F9;
        15'h0CC5: data = 12'h800;
        15'h0CC6: data = 12'h801;
        15'h0CC7: data = 12'h7FF;
        15'h0CC8: data = 12'h803;
        15'h0CC9: data = 12'h7FF;
        15'h0CCA: data = 12'h7F8;
        15'h0CCB: data = 12'h7F7;
        15'h0CCC: data = 12'h7F6;
        15'h0CCD: data = 12'h7F9;
        15'h0CCE: data = 12'h7FC;
        15'h0CCF: data = 12'h802;
        15'h0CD0: data = 12'h802;
        15'h0CD1: data = 12'h7D3;
        15'h0CD2: data = 12'h553;
        15'h0CD3: data = 12'h069;
        15'h0CD4: data = 12'h653;
        15'h0CD5: data = 12'h6C0;
        15'h0CD6: data = 12'h052;
        15'h0CD7: data = 12'h3D5;
        15'h0CD8: data = 12'h7BC;
        15'h0CD9: data = 12'h1A9;
        15'h0CDA: data = 12'h1C4;
        15'h0CDB: data = 12'h80C;
        15'h0CDC: data = 12'h480;
        15'h0CDD: data = 12'h091;
        15'h0CDE: data = 12'h711;
        15'h0CDF: data = 12'h670;
        15'h0CE0: data = 12'h03E;
        15'h0CE1: data = 12'h423;
        15'h0CE2: data = 12'h7BA;
        15'h0CE3: data = 12'h189;
        15'h0CE4: data = 12'h1D3;
        15'h0CE5: data = 12'h80B;
        15'h0CE6: data = 12'h43E;
        15'h0CE7: data = 12'h09B;
        15'h0CE8: data = 12'h73A;
        15'h0CE9: data = 12'h646;
        15'h0CEA: data = 12'h042;
        15'h0CEB: data = 12'h4DC;
        15'h0CEC: data = 12'h785;
        15'h0CED: data = 12'h0F5;
        15'h0CEE: data = 12'h285;
        15'h0CEF: data = 12'h801;
        15'h0CF0: data = 12'h31B;
        15'h0CF1: data = 12'h0FE;
        15'h0CF2: data = 12'h7AE;
        15'h0CF3: data = 12'h54B;
        15'h0CF4: data = 12'h05B;
        15'h0CF5: data = 12'h5A9;
        15'h0CF6: data = 12'h736;
        15'h0CF7: data = 12'h0BF;
        15'h0CF8: data = 12'h2C9;
        15'h0CF9: data = 12'h7FC;
        15'h0CFA: data = 12'h2EC;
        15'h0CFB: data = 12'h10C;
        15'h0CFC: data = 12'h7BF;
        15'h0CFD: data = 12'h57D;
        15'h0CFE: data = 12'h054;
        15'h0CFF: data = 12'h5C6;
        15'h0D00: data = 12'h738;
        15'h0D01: data = 12'h0AF;
        15'h0D02: data = 12'h321;
        15'h0D03: data = 12'h7F9;
        15'h0D04: data = 12'h2EE;
        15'h0D05: data = 12'h126;
        15'h0D06: data = 12'h7BD;
        15'h0D07: data = 12'h583;
        15'h0D08: data = 12'h05B;
        15'h0D09: data = 12'h5FB;
        15'h0D0A: data = 12'h728;
        15'h0D0B: data = 12'h081;
        15'h0D0C: data = 12'h318;
        15'h0D0D: data = 12'h7F0;
        15'h0D0E: data = 12'h2A8;
        15'h0D0F: data = 12'h14F;
        15'h0D10: data = 12'h7C7;
        15'h0D11: data = 12'h55D;
        15'h0D12: data = 12'h05E;
        15'h0D13: data = 12'h5FF;
        15'h0D14: data = 12'h700;
        15'h0D15: data = 12'h063;
        15'h0D16: data = 12'h37E;
        15'h0D17: data = 12'h7E2;
        15'h0D18: data = 12'h221;
        15'h0D19: data = 12'h17C;
        15'h0D1A: data = 12'h7E4;
        15'h0D1B: data = 12'h4E5;
        15'h0D1C: data = 12'h081;
        15'h0D1D: data = 12'h684;
        15'h0D1E: data = 12'h6A6;
        15'h0D1F: data = 12'h040;
        15'h0D20: data = 12'h40E;
        15'h0D21: data = 12'h7BB;
        15'h0D22: data = 12'h18B;
        15'h0D23: data = 12'h1C8;
        15'h0D24: data = 12'h7FC;
        15'h0D25: data = 12'h3F8;
        15'h0D26: data = 12'h0B6;
        15'h0D27: data = 12'h746;
        15'h0D28: data = 12'h620;
        15'h0D29: data = 12'h03E;
        15'h0D2A: data = 12'h4A7;
        15'h0D2B: data = 12'h798;
        15'h0D2C: data = 12'h146;
        15'h0D2D: data = 12'h25D;
        15'h0D2E: data = 12'h80D;
        15'h0D2F: data = 12'h22A;
        15'h0D30: data = 12'h19B;
        15'h0D31: data = 12'h813;
        15'h0D32: data = 12'h2FB;
        15'h0D33: data = 12'h126;
        15'h0D34: data = 12'h7D2;
        15'h0D35: data = 12'h3E3;
        15'h0D36: data = 12'h0D3;
        15'h0D37: data = 12'h777;
        15'h0D38: data = 12'h4A0;
        15'h0D39: data = 12'h097;
        15'h0D3A: data = 12'h71F;
        15'h0D3B: data = 12'h4E2;
        15'h0D3C: data = 12'h083;
        15'h0D3D: data = 12'h718;
        15'h0D3E: data = 12'h534;
        15'h0D3F: data = 12'h079;
        15'h0D40: data = 12'h6C8;
        15'h0D41: data = 12'h57C;
        15'h0D42: data = 12'h064;
        15'h0D43: data = 12'h5DA;
        15'h0D44: data = 12'h65A;
        15'h0D45: data = 12'h058;
        15'h0D46: data = 12'h523;
        15'h0D47: data = 12'h6B9;
        15'h0D48: data = 12'h055;
        15'h0D49: data = 12'h476;
        15'h0D4A: data = 12'h73D;
        15'h0D4B: data = 12'h0A4;
        15'h0D4C: data = 12'h2F5;
        15'h0D4D: data = 12'h7E1;
        15'h0D4E: data = 12'h1B5;
        15'h0D4F: data = 12'h20E;
        15'h0D50: data = 12'h7EE;
        15'h0D51: data = 12'h1D0;
        15'h0D52: data = 12'h1DF;
        15'h0D53: data = 12'h814;
        15'h0D54: data = 12'h2C4;
        15'h0D55: data = 12'h138;
        15'h0D56: data = 12'h820;
        15'h0D57: data = 12'h2F4;
        15'h0D58: data = 12'h128;
        15'h0D59: data = 12'h821;
        15'h0D5A: data = 12'h36E;
        15'h0D5B: data = 12'h0F2;
        15'h0D5C: data = 12'h7ED;
        15'h0D5D: data = 12'h489;
        15'h0D5E: data = 12'h0A6;
        15'h0D5F: data = 12'h7AE;
        15'h0D60: data = 12'h4EF;
        15'h0D61: data = 12'h085;
        15'h0D62: data = 12'h7A1;
        15'h0D63: data = 12'h47C;
        15'h0D64: data = 12'h0AA;
        15'h0D65: data = 12'h7A9;
        15'h0D66: data = 12'h474;
        15'h0D67: data = 12'h0A1;
        15'h0D68: data = 12'h785;
        15'h0D69: data = 12'h4D4;
        15'h0D6A: data = 12'h081;
        15'h0D6B: data = 12'h74D;
        15'h0D6C: data = 12'h4AF;
        15'h0D6D: data = 12'h089;
        15'h0D6E: data = 12'h077;
        15'h0D6F: data = 12'h07A;
        15'h0D70: data = 12'h07B;
        15'h0D71: data = 12'h07B;
        15'h0D72: data = 12'h07F;
        15'h0D73: data = 12'h07A;
        15'h0D74: data = 12'h080;
        15'h0D75: data = 12'h084;
        15'h0D76: data = 12'h082;
        15'h0D77: data = 12'h085;
        15'h0D78: data = 12'h087;
        15'h0D79: data = 12'h08A;
        15'h0D7A: data = 12'h08D;
        15'h0D7B: data = 12'h08A;
        15'h0D7C: data = 12'h08B;
        15'h0D7D: data = 12'h089;
        15'h0D7E: data = 12'h085;
        15'h0D7F: data = 12'h085;
        15'h0D80: data = 12'h080;
        15'h0D81: data = 12'h081;
        15'h0D82: data = 12'h07F;
        15'h0D83: data = 12'h080;
        15'h0D84: data = 12'h07D;
        15'h0D85: data = 12'h07E;
        15'h0D86: data = 12'h07F;
        15'h0D87: data = 12'h083;
        15'h0D88: data = 12'h089;
        15'h0D89: data = 12'h08A;
        15'h0D8A: data = 12'h08D;
        15'h0D8B: data = 12'h08D;
        15'h0D8C: data = 12'h08F;
        15'h0D8D: data = 12'h091;
        15'h0D8E: data = 12'h088;
        15'h0D8F: data = 12'h087;
        15'h0D90: data = 12'h081;
        15'h0D91: data = 12'h07E;
        15'h0D92: data = 12'h07E;
        15'h0D93: data = 12'h081;
        15'h0D94: data = 12'h087;
        15'h0D95: data = 12'h08D;
        15'h0D96: data = 12'h08C;
        15'h0D97: data = 12'h089;
        15'h0D98: data = 12'h089;
        15'h0D99: data = 12'h08B;
        15'h0D9A: data = 12'h087;
        15'h0D9B: data = 12'h083;
        15'h0D9C: data = 12'h080;
        15'h0D9D: data = 12'h07E;
        15'h0D9E: data = 12'h07E;
        15'h0D9F: data = 12'h082;
        15'h0DA0: data = 12'h089;
        15'h0DA1: data = 12'h08D;
        15'h0DA2: data = 12'h08B;
        15'h0DA3: data = 12'h08B;
        15'h0DA4: data = 12'h085;
        15'h0DA5: data = 12'h07E;
        15'h0DA6: data = 12'h07A;
        15'h0DA7: data = 12'h07B;
        15'h0DA8: data = 12'h07A;
        15'h0DA9: data = 12'h082;
        15'h0DAA: data = 12'h086;
        15'h0DAB: data = 12'h08C;
        15'h0DAC: data = 12'h08C;
        15'h0DAD: data = 12'h089;
        15'h0DAE: data = 12'h081;
        15'h0DAF: data = 12'h081;
        15'h0DB0: data = 12'h09D;
        15'h0DB1: data = 12'h0A0;
        15'h0DB2: data = 12'h0A3;
        15'h0DB3: data = 12'h0A8;
        15'h0DB4: data = 12'h0AB;
        15'h0DB5: data = 12'h0AD;
        15'h0DB6: data = 12'h0AB;
        15'h0DB7: data = 12'h0A7;
        15'h0DB8: data = 12'h0A0;
        15'h0DB9: data = 12'h09B;
        15'h0DBA: data = 12'h0A1;
        15'h0DBB: data = 12'h0A5;
        15'h0DBC: data = 12'h0A9;
        15'h0DBD: data = 12'h0AD;
        15'h0DBE: data = 12'h0AC;
        15'h0DBF: data = 12'h0A8;
        15'h0DC0: data = 12'h0A3;
        15'h0DC1: data = 12'h09C;
        15'h0DC2: data = 12'h09A;
        15'h0DC3: data = 12'h09B;
        15'h0DC4: data = 12'h0A3;
        15'h0DC5: data = 12'h0A7;
        15'h0DC6: data = 12'h0A9;
        15'h0DC7: data = 12'h0A9;
        15'h0DC8: data = 12'h0A8;
        15'h0DC9: data = 12'h0A3;
        15'h0DCA: data = 12'h09F;
        15'h0DCB: data = 12'h09F;
        15'h0DCC: data = 12'h09E;
        15'h0DCD: data = 12'h0A1;
        15'h0DCE: data = 12'h0A5;
        15'h0DCF: data = 12'h0AD;
        15'h0DD0: data = 12'h0AD;
        15'h0DD1: data = 12'h0A7;
        15'h0DD2: data = 12'h0A3;
        15'h0DD3: data = 12'h09A;
        15'h0DD4: data = 12'h09A;
        15'h0DD5: data = 12'h09C;
        15'h0DD6: data = 12'h0A3;
        15'h0DD7: data = 12'h0A9;
        15'h0DD8: data = 12'h0AA;
        15'h0DD9: data = 12'h0AB;
        15'h0DDA: data = 12'h0A5;
        15'h0DDB: data = 12'h0A5;
        15'h0DDC: data = 12'h0A2;
        15'h0DDD: data = 12'h0A1;
        15'h0DDE: data = 12'h09E;
        15'h0DDF: data = 12'h09C;
        15'h0DE0: data = 12'h0A4;
        15'h0DE1: data = 12'h0A5;
        15'h0DE2: data = 12'h0AB;
        15'h0DE3: data = 12'h0AB;
        15'h0DE4: data = 12'h0A7;
        15'h0DE5: data = 12'h0A3;
        15'h0DE6: data = 12'h0A1;
        15'h0DE7: data = 12'h09C;
        15'h0DE8: data = 12'h09D;
        15'h0DE9: data = 12'h09A;
        15'h0DEA: data = 12'h0A4;
        15'h0DEB: data = 12'h0AA;
        15'h0DEC: data = 12'h0A9;
        15'h0DED: data = 12'h0AA;
        15'h0DEE: data = 12'h0A8;
        15'h0DEF: data = 12'h0A1;
        15'h0DF0: data = 12'h09C;
        15'h0DF1: data = 12'h09D;
        15'h0DF2: data = 12'h09C;
        15'h0DF3: data = 12'h09C;
        15'h0DF4: data = 12'h0A5;
        15'h0DF5: data = 12'h0A9;
        15'h0DF6: data = 12'h0A9;
        15'h0DF7: data = 12'h0A9;
        15'h0DF8: data = 12'h0A3;
        15'h0DF9: data = 12'h0A4;
        15'h0DFA: data = 12'h0A1;
        15'h0DFB: data = 12'h09F;
        15'h0DFC: data = 12'h09C;
        15'h0DFD: data = 12'h09F;
        15'h0DFE: data = 12'h0BD;
        15'h0DFF: data = 12'h0C5;
        15'h0E00: data = 12'h0C7;
        15'h0E01: data = 12'h0C6;
        15'h0E02: data = 12'h0C6;
        15'h0E03: data = 12'h0C5;
        15'h0E04: data = 12'h0C5;
        15'h0E05: data = 12'h0C5;
        15'h0E06: data = 12'h0BE;
        15'h0E07: data = 12'h0C0;
        15'h0E08: data = 12'h0BC;
        15'h0E09: data = 12'h0BF;
        15'h0E0A: data = 12'h0C0;
        15'h0E0B: data = 12'h0C3;
        15'h0E0C: data = 12'h0C6;
        15'h0E0D: data = 12'h0CA;
        15'h0E0E: data = 12'h0CE;
        15'h0E0F: data = 12'h0C7;
        15'h0E10: data = 12'h0C7;
        15'h0E11: data = 12'h0BD;
        15'h0E12: data = 12'h0BB;
        15'h0E13: data = 12'h0BB;
        15'h0E14: data = 12'h0BD;
        15'h0E15: data = 12'h0BF;
        15'h0E16: data = 12'h0C5;
        15'h0E17: data = 12'h0C6;
        15'h0E18: data = 12'h0C7;
        15'h0E19: data = 12'h0CB;
        15'h0E1A: data = 12'h0C9;
        15'h0E1B: data = 12'h0C8;
        15'h0E1C: data = 12'h0C3;
        15'h0E1D: data = 12'h0C2;
        15'h0E1E: data = 12'h0BE;
        15'h0E1F: data = 12'h0BD;
        15'h0E20: data = 12'h0BD;
        15'h0E21: data = 12'h0BB;
        15'h0E22: data = 12'h0C0;
        15'h0E23: data = 12'h0C4;
        15'h0E24: data = 12'h0C8;
        15'h0E25: data = 12'h0CB;
        15'h0E26: data = 12'h0C8;
        15'h0E27: data = 12'h0C8;
        15'h0E28: data = 12'h0C6;
        15'h0E29: data = 12'h0BF;
        15'h0E2A: data = 12'h0BE;
        15'h0E2B: data = 12'h0BE;
        15'h0E2C: data = 12'h0BC;
        15'h0E2D: data = 12'h0C0;
        15'h0E2E: data = 12'h0C7;
        15'h0E2F: data = 12'h0C7;
        15'h0E30: data = 12'h0CA;
        15'h0E31: data = 12'h0CB;
        15'h0E32: data = 12'h0CA;
        15'h0E33: data = 12'h0C7;
        15'h0E34: data = 12'h0CA;
        15'h0E35: data = 12'h0C2;
        15'h0E36: data = 12'h0BC;
        15'h0E37: data = 12'h0B9;
        15'h0E38: data = 12'h0BD;
        15'h0E39: data = 12'h0BC;
        15'h0E3A: data = 12'h0BE;
        15'h0E3B: data = 12'h0C1;
        15'h0E3C: data = 12'h0C8;
        15'h0E3D: data = 12'h0CB;
        15'h0E3E: data = 12'h0C8;
        15'h0E3F: data = 12'h0C5;
        15'h0E40: data = 12'h0E8;
        15'h0E41: data = 12'h0E8;
        15'h0E42: data = 12'h0E3;
        15'h0E43: data = 12'h0DF;
        15'h0E44: data = 12'h0E1;
        15'h0E45: data = 12'h0E2;
        15'h0E46: data = 12'h0E1;
        15'h0E47: data = 12'h0E6;
        15'h0E48: data = 12'h0E3;
        15'h0E49: data = 12'h0EA;
        15'h0E4A: data = 12'h0E7;
        15'h0E4B: data = 12'h0E7;
        15'h0E4C: data = 12'h0E8;
        15'h0E4D: data = 12'h0E8;
        15'h0E4E: data = 12'h0E5;
        15'h0E4F: data = 12'h0E0;
        15'h0E50: data = 12'h0DD;
        15'h0E51: data = 12'h0DA;
        15'h0E52: data = 12'h0DB;
        15'h0E53: data = 12'h0E3;
        15'h0E54: data = 12'h0E5;
        15'h0E55: data = 12'h0EB;
        15'h0E56: data = 12'h0E7;
        15'h0E57: data = 12'h0EC;
        15'h0E58: data = 12'h0ED;
        15'h0E59: data = 12'h0E7;
        15'h0E5A: data = 12'h0E2;
        15'h0E5B: data = 12'h0DE;
        15'h0E5C: data = 12'h0E1;
        15'h0E5D: data = 12'h0E0;
        15'h0E5E: data = 12'h0E2;
        15'h0E5F: data = 12'h0E1;
        15'h0E60: data = 12'h0E6;
        15'h0E61: data = 12'h0EB;
        15'h0E62: data = 12'h0EA;
        15'h0E63: data = 12'h0EC;
        15'h0E64: data = 12'h0EB;
        15'h0E65: data = 12'h0E4;
        15'h0E66: data = 12'h0E3;
        15'h0E67: data = 12'h0E0;
        15'h0E68: data = 12'h0DB;
        15'h0E69: data = 12'h0DE;
        15'h0E6A: data = 12'h0DF;
        15'h0E6B: data = 12'h0E5;
        15'h0E6C: data = 12'h0E3;
        15'h0E6D: data = 12'h0E9;
        15'h0E6E: data = 12'h0E8;
        15'h0E6F: data = 12'h0E8;
        15'h0E70: data = 12'h0E8;
        15'h0E71: data = 12'h0E9;
        15'h0E72: data = 12'h0E5;
        15'h0E73: data = 12'h0E0;
        15'h0E74: data = 12'h0DE;
        15'h0E75: data = 12'h0DC;
        15'h0E76: data = 12'h0E3;
        15'h0E77: data = 12'h0E5;
        15'h0E78: data = 12'h0E7;
        15'h0E79: data = 12'h0E9;
        15'h0E7A: data = 12'h0EC;
        15'h0E7B: data = 12'h0EC;
        15'h0E7C: data = 12'h0E4;
        15'h0E7D: data = 12'h0E2;
        15'h0E7E: data = 12'h0E1;
        15'h0E7F: data = 12'h0DE;
        15'h0E80: data = 12'h0DE;
        15'h0E81: data = 12'h0E1;
        15'h0E82: data = 12'h0E1;
        15'h0E83: data = 12'h0E7;
        15'h0E84: data = 12'h0EA;
        15'h0E85: data = 12'h0E9;
        15'h0E86: data = 12'h0E8;
        15'h0E87: data = 12'h0E9;
        15'h0E88: data = 12'h0E7;
        15'h0E89: data = 12'h0E3;
        15'h0E8A: data = 12'h0E4;
        15'h0E8B: data = 12'h0DD;
        15'h0E8C: data = 12'h0DC;
        15'h0E8D: data = 12'h0D9;
        15'h0E8E: data = 12'h0DF;
        15'h0E8F: data = 12'h0E7;
        15'h0E90: data = 12'h0EB;
        15'h0E91: data = 12'h0EC;
        15'h0E92: data = 12'h0EC;
        15'h0E93: data = 12'h0E7;
        15'h0E94: data = 12'h0E4;
        15'h0E95: data = 12'h0DD;
        15'h0E96: data = 12'h0DC;
        15'h0E97: data = 12'h0DE;
        15'h0E98: data = 12'h0DF;
        15'h0E99: data = 12'h0E4;
        15'h0E9A: data = 12'h0E7;
        15'h0E9B: data = 12'h100;
        15'h0E9C: data = 12'h10B;
        15'h0E9D: data = 12'h102;
        15'h0E9E: data = 12'h108;
        15'h0E9F: data = 12'h105;
        15'h0EA0: data = 12'h103;
        15'h0EA1: data = 12'h0FD;
        15'h0EA2: data = 12'h0FF;
        15'h0EA3: data = 12'h0FD;
        15'h0EA4: data = 12'h102;
        15'h0EA5: data = 12'h107;
        15'h0EA6: data = 12'h109;
        15'h0EA7: data = 12'h10A;
        15'h0EA8: data = 12'h109;
        15'h0EA9: data = 12'h108;
        15'h0EAA: data = 12'h108;
        15'h0EAB: data = 12'h102;
        15'h0EAC: data = 12'h102;
        15'h0EAD: data = 12'h103;
        15'h0EAE: data = 12'h0FD;
        15'h0EAF: data = 12'h101;
        15'h0EB0: data = 12'h103;
        15'h0EB1: data = 12'h106;
        15'h0EB2: data = 12'h109;
        15'h0EB3: data = 12'h109;
        15'h0EB4: data = 12'h10B;
        15'h0EB5: data = 12'h106;
        15'h0EB6: data = 12'h102;
        15'h0EB7: data = 12'h0FA;
        15'h0EB8: data = 12'h0FA;
        15'h0EB9: data = 12'h0FE;
        15'h0EBA: data = 12'h101;
        15'h0EBB: data = 12'h103;
        15'h0EBC: data = 12'h108;
        15'h0EBD: data = 12'h109;
        15'h0EBE: data = 12'h106;
        15'h0EBF: data = 12'h108;
        15'h0EC0: data = 12'h108;
        15'h0EC1: data = 12'h108;
        15'h0EC2: data = 12'h105;
        15'h0EC3: data = 12'h102;
        15'h0EC4: data = 12'h0FE;
        15'h0EC5: data = 12'h0FE;
        15'h0EC6: data = 12'h0FF;
        15'h0EC7: data = 12'h105;
        15'h0EC8: data = 12'h108;
        15'h0EC9: data = 12'h10C;
        15'h0ECA: data = 12'h10D;
        15'h0ECB: data = 12'h106;
        15'h0ECC: data = 12'h106;
        15'h0ECD: data = 12'h0FF;
        15'h0ECE: data = 12'h0FF;
        15'h0ECF: data = 12'h0FE;
        15'h0ED0: data = 12'h0FE;
        15'h0ED1: data = 12'h0FE;
        15'h0ED2: data = 12'h104;
        15'h0ED3: data = 12'h109;
        15'h0ED4: data = 12'h10A;
        15'h0ED5: data = 12'h10A;
        15'h0ED6: data = 12'h10B;
        15'h0ED7: data = 12'h109;
        15'h0ED8: data = 12'h104;
        15'h0ED9: data = 12'h102;
        15'h0EDA: data = 12'h0FF;
        15'h0EDB: data = 12'h0FB;
        15'h0EDC: data = 12'h102;
        15'h0EDD: data = 12'h126;
        15'h0EDE: data = 12'h12A;
        15'h0EDF: data = 12'h130;
        15'h0EE0: data = 12'h12D;
        15'h0EE1: data = 12'h130;
        15'h0EE2: data = 12'h12D;
        15'h0EE3: data = 12'h12A;
        15'h0EE4: data = 12'h124;
        15'h0EE5: data = 12'h122;
        15'h0EE6: data = 12'h120;
        15'h0EE7: data = 12'h122;
        15'h0EE8: data = 12'h127;
        15'h0EE9: data = 12'h126;
        15'h0EEA: data = 12'h12B;
        15'h0EEB: data = 12'h12A;
        15'h0EEC: data = 12'h128;
        15'h0EED: data = 12'h12A;
        15'h0EEE: data = 12'h12D;
        15'h0EEF: data = 12'h129;
        15'h0EF0: data = 12'h125;
        15'h0EF1: data = 12'h11D;
        15'h0EF2: data = 12'h11D;
        15'h0EF3: data = 12'h11F;
        15'h0EF4: data = 12'h123;
        15'h0EF5: data = 12'h129;
        15'h0EF6: data = 12'h12C;
        15'h0EF7: data = 12'h12F;
        15'h0EF8: data = 12'h12D;
        15'h0EF9: data = 12'h128;
        15'h0EFA: data = 12'h129;
        15'h0EFB: data = 12'h120;
        15'h0EFC: data = 12'h11C;
        15'h0EFD: data = 12'h11D;
        15'h0EFE: data = 12'h11C;
        15'h0EFF: data = 12'h122;
        15'h0F00: data = 12'h127;
        15'h0F01: data = 12'h12B;
        15'h0F02: data = 12'h12E;
        15'h0F03: data = 12'h12A;
        15'h0F04: data = 12'h127;
        15'h0F05: data = 12'h125;
        15'h0F06: data = 12'h122;
        15'h0F07: data = 12'h121;
        15'h0F08: data = 12'h127;
        15'h0F09: data = 12'h11F;
        15'h0F0A: data = 12'h123;
        15'h0F0B: data = 12'h126;
        15'h0F0C: data = 12'h127;
        15'h0F0D: data = 12'h12A;
        15'h0F0E: data = 12'h128;
        15'h0F0F: data = 12'h12A;
        15'h0F10: data = 12'h12B;
        15'h0F11: data = 12'h128;
        15'h0F12: data = 12'h129;
        15'h0F13: data = 12'h122;
        15'h0F14: data = 12'h11F;
        15'h0F15: data = 12'h11C;
        15'h0F16: data = 12'h11D;
        15'h0F17: data = 12'h122;
        15'h0F18: data = 12'h123;
        15'h0F19: data = 12'h12C;
        15'h0F1A: data = 12'h129;
        15'h0F1B: data = 12'h128;
        15'h0F1C: data = 12'h12A;
        15'h0F1D: data = 12'h126;
        15'h0F1E: data = 12'h123;
        15'h0F1F: data = 12'h133;
        15'h0F20: data = 12'h132;
        15'h0F21: data = 12'h135;
        15'h0F22: data = 12'h134;
        15'h0F23: data = 12'h138;
        15'h0F24: data = 12'h13E;
        15'h0F25: data = 12'h13D;
        15'h0F26: data = 12'h13F;
        15'h0F27: data = 12'h13D;
        15'h0F28: data = 12'h13C;
        15'h0F29: data = 12'h136;
        15'h0F2A: data = 12'h131;
        15'h0F2B: data = 12'h12F;
        15'h0F2C: data = 12'h132;
        15'h0F2D: data = 12'h134;
        15'h0F2E: data = 12'h136;
        15'h0F2F: data = 12'h139;
        15'h0F30: data = 12'h140;
        15'h0F31: data = 12'h13D;
        15'h0F32: data = 12'h143;
        15'h0F33: data = 12'h13D;
        15'h0F34: data = 12'h13B;
        15'h0F35: data = 12'h133;
        15'h0F36: data = 12'h130;
        15'h0F37: data = 12'h132;
        15'h0F38: data = 12'h130;
        15'h0F39: data = 12'h132;
        15'h0F3A: data = 12'h135;
        15'h0F3B: data = 12'h13D;
        15'h0F3C: data = 12'h13C;
        15'h0F3D: data = 12'h141;
        15'h0F3E: data = 12'h13C;
        15'h0F3F: data = 12'h139;
        15'h0F40: data = 12'h13A;
        15'h0F41: data = 12'h134;
        15'h0F42: data = 12'h132;
        15'h0F43: data = 12'h137;
        15'h0F44: data = 12'h135;
        15'h0F45: data = 12'h137;
        15'h0F46: data = 12'h13A;
        15'h0F47: data = 12'h13D;
        15'h0F48: data = 12'h138;
        15'h0F49: data = 12'h139;
        15'h0F4A: data = 12'h13A;
        15'h0F4B: data = 12'h139;
        15'h0F4C: data = 12'h137;
        15'h0F4D: data = 12'h134;
        15'h0F4E: data = 12'h130;
        15'h0F4F: data = 12'h134;
        15'h0F50: data = 12'h134;
        15'h0F51: data = 12'h13B;
        15'h0F52: data = 12'h13D;
        15'h0F53: data = 12'h13F;
        15'h0F54: data = 12'h145;
        default: data = 12'h000;
    endcase
end

endmodule
